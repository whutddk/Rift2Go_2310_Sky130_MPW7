magic
tech sky130A
magscale 1 2
timestamp 1669249183
<< obsli1 >>
rect 1104 2159 540408 649009
<< obsm1 >>
rect 474 2128 541498 649324
<< metal2 >>
rect 8298 650726 8354 651526
rect 23294 650726 23350 651526
rect 38290 650726 38346 651526
rect 53286 650726 53342 651526
rect 68282 650726 68338 651526
rect 83278 650726 83334 651526
rect 98274 650726 98330 651526
rect 113270 650726 113326 651526
rect 128266 650726 128322 651526
rect 143262 650726 143318 651526
rect 158258 650726 158314 651526
rect 173254 650726 173310 651526
rect 188250 650726 188306 651526
rect 203246 650726 203302 651526
rect 218242 650726 218298 651526
rect 233238 650726 233294 651526
rect 248234 650726 248290 651526
rect 263230 650726 263286 651526
rect 278226 650726 278282 651526
rect 293222 650726 293278 651526
rect 308218 650726 308274 651526
rect 323214 650726 323270 651526
rect 338210 650726 338266 651526
rect 353206 650726 353262 651526
rect 368202 650726 368258 651526
rect 383198 650726 383254 651526
rect 398194 650726 398250 651526
rect 413190 650726 413246 651526
rect 428186 650726 428242 651526
rect 443182 650726 443238 651526
rect 458178 650726 458234 651526
rect 473174 650726 473230 651526
rect 488170 650726 488226 651526
rect 503166 650726 503222 651526
rect 518162 650726 518218 651526
rect 533158 650726 533214 651526
rect 21270 0 21326 800
rect 22282 0 22338 800
rect 23294 0 23350 800
rect 24306 0 24362 800
rect 25318 0 25374 800
rect 26330 0 26386 800
rect 27342 0 27398 800
rect 28354 0 28410 800
rect 29366 0 29422 800
rect 30378 0 30434 800
rect 31390 0 31446 800
rect 32402 0 32458 800
rect 33414 0 33470 800
rect 34426 0 34482 800
rect 35438 0 35494 800
rect 36450 0 36506 800
rect 37462 0 37518 800
rect 38474 0 38530 800
rect 39486 0 39542 800
rect 40498 0 40554 800
rect 41510 0 41566 800
rect 42522 0 42578 800
rect 43534 0 43590 800
rect 44546 0 44602 800
rect 45558 0 45614 800
rect 46570 0 46626 800
rect 47582 0 47638 800
rect 48594 0 48650 800
rect 49606 0 49662 800
rect 50618 0 50674 800
rect 51630 0 51686 800
rect 52642 0 52698 800
rect 53654 0 53710 800
rect 54666 0 54722 800
rect 55678 0 55734 800
rect 56690 0 56746 800
rect 57702 0 57758 800
rect 58714 0 58770 800
rect 59726 0 59782 800
rect 60738 0 60794 800
rect 61750 0 61806 800
rect 62762 0 62818 800
rect 63774 0 63830 800
rect 64786 0 64842 800
rect 65798 0 65854 800
rect 66810 0 66866 800
rect 67822 0 67878 800
rect 68834 0 68890 800
rect 69846 0 69902 800
rect 70858 0 70914 800
rect 71870 0 71926 800
rect 72882 0 72938 800
rect 73894 0 73950 800
rect 74906 0 74962 800
rect 75918 0 75974 800
rect 76930 0 76986 800
rect 77942 0 77998 800
rect 78954 0 79010 800
rect 79966 0 80022 800
rect 80978 0 81034 800
rect 81990 0 82046 800
rect 83002 0 83058 800
rect 84014 0 84070 800
rect 85026 0 85082 800
rect 86038 0 86094 800
rect 87050 0 87106 800
rect 88062 0 88118 800
rect 89074 0 89130 800
rect 90086 0 90142 800
rect 91098 0 91154 800
rect 92110 0 92166 800
rect 93122 0 93178 800
rect 94134 0 94190 800
rect 95146 0 95202 800
rect 96158 0 96214 800
rect 97170 0 97226 800
rect 98182 0 98238 800
rect 99194 0 99250 800
rect 100206 0 100262 800
rect 101218 0 101274 800
rect 102230 0 102286 800
rect 103242 0 103298 800
rect 104254 0 104310 800
rect 105266 0 105322 800
rect 106278 0 106334 800
rect 107290 0 107346 800
rect 108302 0 108358 800
rect 109314 0 109370 800
rect 110326 0 110382 800
rect 111338 0 111394 800
rect 112350 0 112406 800
rect 113362 0 113418 800
rect 114374 0 114430 800
rect 115386 0 115442 800
rect 116398 0 116454 800
rect 117410 0 117466 800
rect 118422 0 118478 800
rect 119434 0 119490 800
rect 120446 0 120502 800
rect 121458 0 121514 800
rect 122470 0 122526 800
rect 123482 0 123538 800
rect 124494 0 124550 800
rect 125506 0 125562 800
rect 126518 0 126574 800
rect 127530 0 127586 800
rect 128542 0 128598 800
rect 129554 0 129610 800
rect 130566 0 130622 800
rect 131578 0 131634 800
rect 132590 0 132646 800
rect 133602 0 133658 800
rect 134614 0 134670 800
rect 135626 0 135682 800
rect 136638 0 136694 800
rect 137650 0 137706 800
rect 138662 0 138718 800
rect 139674 0 139730 800
rect 140686 0 140742 800
rect 141698 0 141754 800
rect 142710 0 142766 800
rect 143722 0 143778 800
rect 144734 0 144790 800
rect 145746 0 145802 800
rect 146758 0 146814 800
rect 147770 0 147826 800
rect 148782 0 148838 800
rect 149794 0 149850 800
rect 150806 0 150862 800
rect 151818 0 151874 800
rect 152830 0 152886 800
rect 153842 0 153898 800
rect 154854 0 154910 800
rect 155866 0 155922 800
rect 156878 0 156934 800
rect 157890 0 157946 800
rect 158902 0 158958 800
rect 159914 0 159970 800
rect 160926 0 160982 800
rect 161938 0 161994 800
rect 162950 0 163006 800
rect 163962 0 164018 800
rect 164974 0 165030 800
rect 165986 0 166042 800
rect 166998 0 167054 800
rect 168010 0 168066 800
rect 169022 0 169078 800
rect 170034 0 170090 800
rect 171046 0 171102 800
rect 172058 0 172114 800
rect 173070 0 173126 800
rect 174082 0 174138 800
rect 175094 0 175150 800
rect 176106 0 176162 800
rect 177118 0 177174 800
rect 178130 0 178186 800
rect 179142 0 179198 800
rect 180154 0 180210 800
rect 181166 0 181222 800
rect 182178 0 182234 800
rect 183190 0 183246 800
rect 184202 0 184258 800
rect 185214 0 185270 800
rect 186226 0 186282 800
rect 187238 0 187294 800
rect 188250 0 188306 800
rect 189262 0 189318 800
rect 190274 0 190330 800
rect 191286 0 191342 800
rect 192298 0 192354 800
rect 193310 0 193366 800
rect 194322 0 194378 800
rect 195334 0 195390 800
rect 196346 0 196402 800
rect 197358 0 197414 800
rect 198370 0 198426 800
rect 199382 0 199438 800
rect 200394 0 200450 800
rect 201406 0 201462 800
rect 202418 0 202474 800
rect 203430 0 203486 800
rect 204442 0 204498 800
rect 205454 0 205510 800
rect 206466 0 206522 800
rect 207478 0 207534 800
rect 208490 0 208546 800
rect 209502 0 209558 800
rect 210514 0 210570 800
rect 211526 0 211582 800
rect 212538 0 212594 800
rect 213550 0 213606 800
rect 214562 0 214618 800
rect 215574 0 215630 800
rect 216586 0 216642 800
rect 217598 0 217654 800
rect 218610 0 218666 800
rect 219622 0 219678 800
rect 220634 0 220690 800
rect 221646 0 221702 800
rect 222658 0 222714 800
rect 223670 0 223726 800
rect 224682 0 224738 800
rect 225694 0 225750 800
rect 226706 0 226762 800
rect 227718 0 227774 800
rect 228730 0 228786 800
rect 229742 0 229798 800
rect 230754 0 230810 800
rect 231766 0 231822 800
rect 232778 0 232834 800
rect 233790 0 233846 800
rect 234802 0 234858 800
rect 235814 0 235870 800
rect 236826 0 236882 800
rect 237838 0 237894 800
rect 238850 0 238906 800
rect 239862 0 239918 800
rect 240874 0 240930 800
rect 241886 0 241942 800
rect 242898 0 242954 800
rect 243910 0 243966 800
rect 244922 0 244978 800
rect 245934 0 245990 800
rect 246946 0 247002 800
rect 247958 0 248014 800
rect 248970 0 249026 800
rect 249982 0 250038 800
rect 250994 0 251050 800
rect 252006 0 252062 800
rect 253018 0 253074 800
rect 254030 0 254086 800
rect 255042 0 255098 800
rect 256054 0 256110 800
rect 257066 0 257122 800
rect 258078 0 258134 800
rect 259090 0 259146 800
rect 260102 0 260158 800
rect 261114 0 261170 800
rect 262126 0 262182 800
rect 263138 0 263194 800
rect 264150 0 264206 800
rect 265162 0 265218 800
rect 266174 0 266230 800
rect 267186 0 267242 800
rect 268198 0 268254 800
rect 269210 0 269266 800
rect 270222 0 270278 800
rect 271234 0 271290 800
rect 272246 0 272302 800
rect 273258 0 273314 800
rect 274270 0 274326 800
rect 275282 0 275338 800
rect 276294 0 276350 800
rect 277306 0 277362 800
rect 278318 0 278374 800
rect 279330 0 279386 800
rect 280342 0 280398 800
rect 281354 0 281410 800
rect 282366 0 282422 800
rect 283378 0 283434 800
rect 284390 0 284446 800
rect 285402 0 285458 800
rect 286414 0 286470 800
rect 287426 0 287482 800
rect 288438 0 288494 800
rect 289450 0 289506 800
rect 290462 0 290518 800
rect 291474 0 291530 800
rect 292486 0 292542 800
rect 293498 0 293554 800
rect 294510 0 294566 800
rect 295522 0 295578 800
rect 296534 0 296590 800
rect 297546 0 297602 800
rect 298558 0 298614 800
rect 299570 0 299626 800
rect 300582 0 300638 800
rect 301594 0 301650 800
rect 302606 0 302662 800
rect 303618 0 303674 800
rect 304630 0 304686 800
rect 305642 0 305698 800
rect 306654 0 306710 800
rect 307666 0 307722 800
rect 308678 0 308734 800
rect 309690 0 309746 800
rect 310702 0 310758 800
rect 311714 0 311770 800
rect 312726 0 312782 800
rect 313738 0 313794 800
rect 314750 0 314806 800
rect 315762 0 315818 800
rect 316774 0 316830 800
rect 317786 0 317842 800
rect 318798 0 318854 800
rect 319810 0 319866 800
rect 320822 0 320878 800
rect 321834 0 321890 800
rect 322846 0 322902 800
rect 323858 0 323914 800
rect 324870 0 324926 800
rect 325882 0 325938 800
rect 326894 0 326950 800
rect 327906 0 327962 800
rect 328918 0 328974 800
rect 329930 0 329986 800
rect 330942 0 330998 800
rect 331954 0 332010 800
rect 332966 0 333022 800
rect 333978 0 334034 800
rect 334990 0 335046 800
rect 336002 0 336058 800
rect 337014 0 337070 800
rect 338026 0 338082 800
rect 339038 0 339094 800
rect 340050 0 340106 800
rect 341062 0 341118 800
rect 342074 0 342130 800
rect 343086 0 343142 800
rect 344098 0 344154 800
rect 345110 0 345166 800
rect 346122 0 346178 800
rect 347134 0 347190 800
rect 348146 0 348202 800
rect 349158 0 349214 800
rect 350170 0 350226 800
rect 351182 0 351238 800
rect 352194 0 352250 800
rect 353206 0 353262 800
rect 354218 0 354274 800
rect 355230 0 355286 800
rect 356242 0 356298 800
rect 357254 0 357310 800
rect 358266 0 358322 800
rect 359278 0 359334 800
rect 360290 0 360346 800
rect 361302 0 361358 800
rect 362314 0 362370 800
rect 363326 0 363382 800
rect 364338 0 364394 800
rect 365350 0 365406 800
rect 366362 0 366418 800
rect 367374 0 367430 800
rect 368386 0 368442 800
rect 369398 0 369454 800
rect 370410 0 370466 800
rect 371422 0 371478 800
rect 372434 0 372490 800
rect 373446 0 373502 800
rect 374458 0 374514 800
rect 375470 0 375526 800
rect 376482 0 376538 800
rect 377494 0 377550 800
rect 378506 0 378562 800
rect 379518 0 379574 800
rect 380530 0 380586 800
rect 381542 0 381598 800
rect 382554 0 382610 800
rect 383566 0 383622 800
rect 384578 0 384634 800
rect 385590 0 385646 800
rect 386602 0 386658 800
rect 387614 0 387670 800
rect 388626 0 388682 800
rect 389638 0 389694 800
rect 390650 0 390706 800
rect 391662 0 391718 800
rect 392674 0 392730 800
rect 393686 0 393742 800
rect 394698 0 394754 800
rect 395710 0 395766 800
rect 396722 0 396778 800
rect 397734 0 397790 800
rect 398746 0 398802 800
rect 399758 0 399814 800
rect 400770 0 400826 800
rect 401782 0 401838 800
rect 402794 0 402850 800
rect 403806 0 403862 800
rect 404818 0 404874 800
rect 405830 0 405886 800
rect 406842 0 406898 800
rect 407854 0 407910 800
rect 408866 0 408922 800
rect 409878 0 409934 800
rect 410890 0 410946 800
rect 411902 0 411958 800
rect 412914 0 412970 800
rect 413926 0 413982 800
rect 414938 0 414994 800
rect 415950 0 416006 800
rect 416962 0 417018 800
rect 417974 0 418030 800
rect 418986 0 419042 800
rect 419998 0 420054 800
rect 421010 0 421066 800
rect 422022 0 422078 800
rect 423034 0 423090 800
rect 424046 0 424102 800
rect 425058 0 425114 800
rect 426070 0 426126 800
rect 427082 0 427138 800
rect 428094 0 428150 800
rect 429106 0 429162 800
rect 430118 0 430174 800
rect 431130 0 431186 800
rect 432142 0 432198 800
rect 433154 0 433210 800
rect 434166 0 434222 800
rect 435178 0 435234 800
rect 436190 0 436246 800
rect 437202 0 437258 800
rect 438214 0 438270 800
rect 439226 0 439282 800
rect 440238 0 440294 800
rect 441250 0 441306 800
rect 442262 0 442318 800
rect 443274 0 443330 800
rect 444286 0 444342 800
rect 445298 0 445354 800
rect 446310 0 446366 800
rect 447322 0 447378 800
rect 448334 0 448390 800
rect 449346 0 449402 800
rect 450358 0 450414 800
rect 451370 0 451426 800
rect 452382 0 452438 800
rect 453394 0 453450 800
rect 454406 0 454462 800
rect 455418 0 455474 800
rect 456430 0 456486 800
rect 457442 0 457498 800
rect 458454 0 458510 800
rect 459466 0 459522 800
rect 460478 0 460534 800
rect 461490 0 461546 800
rect 462502 0 462558 800
rect 463514 0 463570 800
rect 464526 0 464582 800
rect 465538 0 465594 800
rect 466550 0 466606 800
rect 467562 0 467618 800
rect 468574 0 468630 800
rect 469586 0 469642 800
rect 470598 0 470654 800
rect 471610 0 471666 800
rect 472622 0 472678 800
rect 473634 0 473690 800
rect 474646 0 474702 800
rect 475658 0 475714 800
rect 476670 0 476726 800
rect 477682 0 477738 800
rect 478694 0 478750 800
rect 479706 0 479762 800
rect 480718 0 480774 800
rect 481730 0 481786 800
rect 482742 0 482798 800
rect 483754 0 483810 800
rect 484766 0 484822 800
rect 485778 0 485834 800
rect 486790 0 486846 800
rect 487802 0 487858 800
rect 488814 0 488870 800
rect 489826 0 489882 800
rect 490838 0 490894 800
rect 491850 0 491906 800
rect 492862 0 492918 800
rect 493874 0 493930 800
rect 494886 0 494942 800
rect 495898 0 495954 800
rect 496910 0 496966 800
rect 497922 0 497978 800
rect 498934 0 498990 800
rect 499946 0 500002 800
rect 500958 0 501014 800
rect 501970 0 502026 800
rect 502982 0 503038 800
rect 503994 0 504050 800
rect 505006 0 505062 800
rect 506018 0 506074 800
rect 507030 0 507086 800
rect 508042 0 508098 800
rect 509054 0 509110 800
rect 510066 0 510122 800
rect 511078 0 511134 800
rect 512090 0 512146 800
rect 513102 0 513158 800
rect 514114 0 514170 800
rect 515126 0 515182 800
rect 516138 0 516194 800
rect 517150 0 517206 800
rect 518162 0 518218 800
rect 519174 0 519230 800
rect 520186 0 520242 800
<< obsm2 >>
rect 478 650670 8242 650842
rect 8410 650670 23238 650842
rect 23406 650670 38234 650842
rect 38402 650670 53230 650842
rect 53398 650670 68226 650842
rect 68394 650670 83222 650842
rect 83390 650670 98218 650842
rect 98386 650670 113214 650842
rect 113382 650670 128210 650842
rect 128378 650670 143206 650842
rect 143374 650670 158202 650842
rect 158370 650670 173198 650842
rect 173366 650670 188194 650842
rect 188362 650670 203190 650842
rect 203358 650670 218186 650842
rect 218354 650670 233182 650842
rect 233350 650670 248178 650842
rect 248346 650670 263174 650842
rect 263342 650670 278170 650842
rect 278338 650670 293166 650842
rect 293334 650670 308162 650842
rect 308330 650670 323158 650842
rect 323326 650670 338154 650842
rect 338322 650670 353150 650842
rect 353318 650670 368146 650842
rect 368314 650670 383142 650842
rect 383310 650670 398138 650842
rect 398306 650670 413134 650842
rect 413302 650670 428130 650842
rect 428298 650670 443126 650842
rect 443294 650670 458122 650842
rect 458290 650670 473118 650842
rect 473286 650670 488114 650842
rect 488282 650670 503110 650842
rect 503278 650670 518106 650842
rect 518274 650670 533102 650842
rect 533270 650670 541492 650842
rect 478 856 541492 650670
rect 478 734 21214 856
rect 21382 734 22226 856
rect 22394 734 23238 856
rect 23406 734 24250 856
rect 24418 734 25262 856
rect 25430 734 26274 856
rect 26442 734 27286 856
rect 27454 734 28298 856
rect 28466 734 29310 856
rect 29478 734 30322 856
rect 30490 734 31334 856
rect 31502 734 32346 856
rect 32514 734 33358 856
rect 33526 734 34370 856
rect 34538 734 35382 856
rect 35550 734 36394 856
rect 36562 734 37406 856
rect 37574 734 38418 856
rect 38586 734 39430 856
rect 39598 734 40442 856
rect 40610 734 41454 856
rect 41622 734 42466 856
rect 42634 734 43478 856
rect 43646 734 44490 856
rect 44658 734 45502 856
rect 45670 734 46514 856
rect 46682 734 47526 856
rect 47694 734 48538 856
rect 48706 734 49550 856
rect 49718 734 50562 856
rect 50730 734 51574 856
rect 51742 734 52586 856
rect 52754 734 53598 856
rect 53766 734 54610 856
rect 54778 734 55622 856
rect 55790 734 56634 856
rect 56802 734 57646 856
rect 57814 734 58658 856
rect 58826 734 59670 856
rect 59838 734 60682 856
rect 60850 734 61694 856
rect 61862 734 62706 856
rect 62874 734 63718 856
rect 63886 734 64730 856
rect 64898 734 65742 856
rect 65910 734 66754 856
rect 66922 734 67766 856
rect 67934 734 68778 856
rect 68946 734 69790 856
rect 69958 734 70802 856
rect 70970 734 71814 856
rect 71982 734 72826 856
rect 72994 734 73838 856
rect 74006 734 74850 856
rect 75018 734 75862 856
rect 76030 734 76874 856
rect 77042 734 77886 856
rect 78054 734 78898 856
rect 79066 734 79910 856
rect 80078 734 80922 856
rect 81090 734 81934 856
rect 82102 734 82946 856
rect 83114 734 83958 856
rect 84126 734 84970 856
rect 85138 734 85982 856
rect 86150 734 86994 856
rect 87162 734 88006 856
rect 88174 734 89018 856
rect 89186 734 90030 856
rect 90198 734 91042 856
rect 91210 734 92054 856
rect 92222 734 93066 856
rect 93234 734 94078 856
rect 94246 734 95090 856
rect 95258 734 96102 856
rect 96270 734 97114 856
rect 97282 734 98126 856
rect 98294 734 99138 856
rect 99306 734 100150 856
rect 100318 734 101162 856
rect 101330 734 102174 856
rect 102342 734 103186 856
rect 103354 734 104198 856
rect 104366 734 105210 856
rect 105378 734 106222 856
rect 106390 734 107234 856
rect 107402 734 108246 856
rect 108414 734 109258 856
rect 109426 734 110270 856
rect 110438 734 111282 856
rect 111450 734 112294 856
rect 112462 734 113306 856
rect 113474 734 114318 856
rect 114486 734 115330 856
rect 115498 734 116342 856
rect 116510 734 117354 856
rect 117522 734 118366 856
rect 118534 734 119378 856
rect 119546 734 120390 856
rect 120558 734 121402 856
rect 121570 734 122414 856
rect 122582 734 123426 856
rect 123594 734 124438 856
rect 124606 734 125450 856
rect 125618 734 126462 856
rect 126630 734 127474 856
rect 127642 734 128486 856
rect 128654 734 129498 856
rect 129666 734 130510 856
rect 130678 734 131522 856
rect 131690 734 132534 856
rect 132702 734 133546 856
rect 133714 734 134558 856
rect 134726 734 135570 856
rect 135738 734 136582 856
rect 136750 734 137594 856
rect 137762 734 138606 856
rect 138774 734 139618 856
rect 139786 734 140630 856
rect 140798 734 141642 856
rect 141810 734 142654 856
rect 142822 734 143666 856
rect 143834 734 144678 856
rect 144846 734 145690 856
rect 145858 734 146702 856
rect 146870 734 147714 856
rect 147882 734 148726 856
rect 148894 734 149738 856
rect 149906 734 150750 856
rect 150918 734 151762 856
rect 151930 734 152774 856
rect 152942 734 153786 856
rect 153954 734 154798 856
rect 154966 734 155810 856
rect 155978 734 156822 856
rect 156990 734 157834 856
rect 158002 734 158846 856
rect 159014 734 159858 856
rect 160026 734 160870 856
rect 161038 734 161882 856
rect 162050 734 162894 856
rect 163062 734 163906 856
rect 164074 734 164918 856
rect 165086 734 165930 856
rect 166098 734 166942 856
rect 167110 734 167954 856
rect 168122 734 168966 856
rect 169134 734 169978 856
rect 170146 734 170990 856
rect 171158 734 172002 856
rect 172170 734 173014 856
rect 173182 734 174026 856
rect 174194 734 175038 856
rect 175206 734 176050 856
rect 176218 734 177062 856
rect 177230 734 178074 856
rect 178242 734 179086 856
rect 179254 734 180098 856
rect 180266 734 181110 856
rect 181278 734 182122 856
rect 182290 734 183134 856
rect 183302 734 184146 856
rect 184314 734 185158 856
rect 185326 734 186170 856
rect 186338 734 187182 856
rect 187350 734 188194 856
rect 188362 734 189206 856
rect 189374 734 190218 856
rect 190386 734 191230 856
rect 191398 734 192242 856
rect 192410 734 193254 856
rect 193422 734 194266 856
rect 194434 734 195278 856
rect 195446 734 196290 856
rect 196458 734 197302 856
rect 197470 734 198314 856
rect 198482 734 199326 856
rect 199494 734 200338 856
rect 200506 734 201350 856
rect 201518 734 202362 856
rect 202530 734 203374 856
rect 203542 734 204386 856
rect 204554 734 205398 856
rect 205566 734 206410 856
rect 206578 734 207422 856
rect 207590 734 208434 856
rect 208602 734 209446 856
rect 209614 734 210458 856
rect 210626 734 211470 856
rect 211638 734 212482 856
rect 212650 734 213494 856
rect 213662 734 214506 856
rect 214674 734 215518 856
rect 215686 734 216530 856
rect 216698 734 217542 856
rect 217710 734 218554 856
rect 218722 734 219566 856
rect 219734 734 220578 856
rect 220746 734 221590 856
rect 221758 734 222602 856
rect 222770 734 223614 856
rect 223782 734 224626 856
rect 224794 734 225638 856
rect 225806 734 226650 856
rect 226818 734 227662 856
rect 227830 734 228674 856
rect 228842 734 229686 856
rect 229854 734 230698 856
rect 230866 734 231710 856
rect 231878 734 232722 856
rect 232890 734 233734 856
rect 233902 734 234746 856
rect 234914 734 235758 856
rect 235926 734 236770 856
rect 236938 734 237782 856
rect 237950 734 238794 856
rect 238962 734 239806 856
rect 239974 734 240818 856
rect 240986 734 241830 856
rect 241998 734 242842 856
rect 243010 734 243854 856
rect 244022 734 244866 856
rect 245034 734 245878 856
rect 246046 734 246890 856
rect 247058 734 247902 856
rect 248070 734 248914 856
rect 249082 734 249926 856
rect 250094 734 250938 856
rect 251106 734 251950 856
rect 252118 734 252962 856
rect 253130 734 253974 856
rect 254142 734 254986 856
rect 255154 734 255998 856
rect 256166 734 257010 856
rect 257178 734 258022 856
rect 258190 734 259034 856
rect 259202 734 260046 856
rect 260214 734 261058 856
rect 261226 734 262070 856
rect 262238 734 263082 856
rect 263250 734 264094 856
rect 264262 734 265106 856
rect 265274 734 266118 856
rect 266286 734 267130 856
rect 267298 734 268142 856
rect 268310 734 269154 856
rect 269322 734 270166 856
rect 270334 734 271178 856
rect 271346 734 272190 856
rect 272358 734 273202 856
rect 273370 734 274214 856
rect 274382 734 275226 856
rect 275394 734 276238 856
rect 276406 734 277250 856
rect 277418 734 278262 856
rect 278430 734 279274 856
rect 279442 734 280286 856
rect 280454 734 281298 856
rect 281466 734 282310 856
rect 282478 734 283322 856
rect 283490 734 284334 856
rect 284502 734 285346 856
rect 285514 734 286358 856
rect 286526 734 287370 856
rect 287538 734 288382 856
rect 288550 734 289394 856
rect 289562 734 290406 856
rect 290574 734 291418 856
rect 291586 734 292430 856
rect 292598 734 293442 856
rect 293610 734 294454 856
rect 294622 734 295466 856
rect 295634 734 296478 856
rect 296646 734 297490 856
rect 297658 734 298502 856
rect 298670 734 299514 856
rect 299682 734 300526 856
rect 300694 734 301538 856
rect 301706 734 302550 856
rect 302718 734 303562 856
rect 303730 734 304574 856
rect 304742 734 305586 856
rect 305754 734 306598 856
rect 306766 734 307610 856
rect 307778 734 308622 856
rect 308790 734 309634 856
rect 309802 734 310646 856
rect 310814 734 311658 856
rect 311826 734 312670 856
rect 312838 734 313682 856
rect 313850 734 314694 856
rect 314862 734 315706 856
rect 315874 734 316718 856
rect 316886 734 317730 856
rect 317898 734 318742 856
rect 318910 734 319754 856
rect 319922 734 320766 856
rect 320934 734 321778 856
rect 321946 734 322790 856
rect 322958 734 323802 856
rect 323970 734 324814 856
rect 324982 734 325826 856
rect 325994 734 326838 856
rect 327006 734 327850 856
rect 328018 734 328862 856
rect 329030 734 329874 856
rect 330042 734 330886 856
rect 331054 734 331898 856
rect 332066 734 332910 856
rect 333078 734 333922 856
rect 334090 734 334934 856
rect 335102 734 335946 856
rect 336114 734 336958 856
rect 337126 734 337970 856
rect 338138 734 338982 856
rect 339150 734 339994 856
rect 340162 734 341006 856
rect 341174 734 342018 856
rect 342186 734 343030 856
rect 343198 734 344042 856
rect 344210 734 345054 856
rect 345222 734 346066 856
rect 346234 734 347078 856
rect 347246 734 348090 856
rect 348258 734 349102 856
rect 349270 734 350114 856
rect 350282 734 351126 856
rect 351294 734 352138 856
rect 352306 734 353150 856
rect 353318 734 354162 856
rect 354330 734 355174 856
rect 355342 734 356186 856
rect 356354 734 357198 856
rect 357366 734 358210 856
rect 358378 734 359222 856
rect 359390 734 360234 856
rect 360402 734 361246 856
rect 361414 734 362258 856
rect 362426 734 363270 856
rect 363438 734 364282 856
rect 364450 734 365294 856
rect 365462 734 366306 856
rect 366474 734 367318 856
rect 367486 734 368330 856
rect 368498 734 369342 856
rect 369510 734 370354 856
rect 370522 734 371366 856
rect 371534 734 372378 856
rect 372546 734 373390 856
rect 373558 734 374402 856
rect 374570 734 375414 856
rect 375582 734 376426 856
rect 376594 734 377438 856
rect 377606 734 378450 856
rect 378618 734 379462 856
rect 379630 734 380474 856
rect 380642 734 381486 856
rect 381654 734 382498 856
rect 382666 734 383510 856
rect 383678 734 384522 856
rect 384690 734 385534 856
rect 385702 734 386546 856
rect 386714 734 387558 856
rect 387726 734 388570 856
rect 388738 734 389582 856
rect 389750 734 390594 856
rect 390762 734 391606 856
rect 391774 734 392618 856
rect 392786 734 393630 856
rect 393798 734 394642 856
rect 394810 734 395654 856
rect 395822 734 396666 856
rect 396834 734 397678 856
rect 397846 734 398690 856
rect 398858 734 399702 856
rect 399870 734 400714 856
rect 400882 734 401726 856
rect 401894 734 402738 856
rect 402906 734 403750 856
rect 403918 734 404762 856
rect 404930 734 405774 856
rect 405942 734 406786 856
rect 406954 734 407798 856
rect 407966 734 408810 856
rect 408978 734 409822 856
rect 409990 734 410834 856
rect 411002 734 411846 856
rect 412014 734 412858 856
rect 413026 734 413870 856
rect 414038 734 414882 856
rect 415050 734 415894 856
rect 416062 734 416906 856
rect 417074 734 417918 856
rect 418086 734 418930 856
rect 419098 734 419942 856
rect 420110 734 420954 856
rect 421122 734 421966 856
rect 422134 734 422978 856
rect 423146 734 423990 856
rect 424158 734 425002 856
rect 425170 734 426014 856
rect 426182 734 427026 856
rect 427194 734 428038 856
rect 428206 734 429050 856
rect 429218 734 430062 856
rect 430230 734 431074 856
rect 431242 734 432086 856
rect 432254 734 433098 856
rect 433266 734 434110 856
rect 434278 734 435122 856
rect 435290 734 436134 856
rect 436302 734 437146 856
rect 437314 734 438158 856
rect 438326 734 439170 856
rect 439338 734 440182 856
rect 440350 734 441194 856
rect 441362 734 442206 856
rect 442374 734 443218 856
rect 443386 734 444230 856
rect 444398 734 445242 856
rect 445410 734 446254 856
rect 446422 734 447266 856
rect 447434 734 448278 856
rect 448446 734 449290 856
rect 449458 734 450302 856
rect 450470 734 451314 856
rect 451482 734 452326 856
rect 452494 734 453338 856
rect 453506 734 454350 856
rect 454518 734 455362 856
rect 455530 734 456374 856
rect 456542 734 457386 856
rect 457554 734 458398 856
rect 458566 734 459410 856
rect 459578 734 460422 856
rect 460590 734 461434 856
rect 461602 734 462446 856
rect 462614 734 463458 856
rect 463626 734 464470 856
rect 464638 734 465482 856
rect 465650 734 466494 856
rect 466662 734 467506 856
rect 467674 734 468518 856
rect 468686 734 469530 856
rect 469698 734 470542 856
rect 470710 734 471554 856
rect 471722 734 472566 856
rect 472734 734 473578 856
rect 473746 734 474590 856
rect 474758 734 475602 856
rect 475770 734 476614 856
rect 476782 734 477626 856
rect 477794 734 478638 856
rect 478806 734 479650 856
rect 479818 734 480662 856
rect 480830 734 481674 856
rect 481842 734 482686 856
rect 482854 734 483698 856
rect 483866 734 484710 856
rect 484878 734 485722 856
rect 485890 734 486734 856
rect 486902 734 487746 856
rect 487914 734 488758 856
rect 488926 734 489770 856
rect 489938 734 490782 856
rect 490950 734 491794 856
rect 491962 734 492806 856
rect 492974 734 493818 856
rect 493986 734 494830 856
rect 494998 734 495842 856
rect 496010 734 496854 856
rect 497022 734 497866 856
rect 498034 734 498878 856
rect 499046 734 499890 856
rect 500058 734 500902 856
rect 501070 734 501914 856
rect 502082 734 502926 856
rect 503094 734 503938 856
rect 504106 734 504950 856
rect 505118 734 505962 856
rect 506130 734 506974 856
rect 507142 734 507986 856
rect 508154 734 508998 856
rect 509166 734 510010 856
rect 510178 734 511022 856
rect 511190 734 512034 856
rect 512202 734 513046 856
rect 513214 734 514058 856
rect 514226 734 515070 856
rect 515238 734 516082 856
rect 516250 734 517094 856
rect 517262 734 518106 856
rect 518274 734 519118 856
rect 519286 734 520130 856
rect 520298 734 541492 856
<< metal3 >>
rect 540720 643832 541520 643952
rect 0 642744 800 642864
rect 540720 631592 541520 631712
rect 0 630776 800 630896
rect 540720 619352 541520 619472
rect 0 618808 800 618928
rect 540720 607112 541520 607232
rect 0 606840 800 606960
rect 0 594872 800 594992
rect 540720 594872 541520 594992
rect 0 582904 800 583024
rect 540720 582632 541520 582752
rect 0 570936 800 571056
rect 540720 570392 541520 570512
rect 0 558968 800 559088
rect 540720 558152 541520 558272
rect 0 547000 800 547120
rect 540720 545912 541520 546032
rect 0 535032 800 535152
rect 540720 533672 541520 533792
rect 0 523064 800 523184
rect 540720 521432 541520 521552
rect 0 511096 800 511216
rect 540720 509192 541520 509312
rect 0 499128 800 499248
rect 540720 496952 541520 497072
rect 0 487160 800 487280
rect 540720 484712 541520 484832
rect 0 475192 800 475312
rect 540720 472472 541520 472592
rect 0 463224 800 463344
rect 540720 460232 541520 460352
rect 0 451256 800 451376
rect 540720 447992 541520 448112
rect 0 439288 800 439408
rect 540720 435752 541520 435872
rect 0 427320 800 427440
rect 540720 423512 541520 423632
rect 0 415352 800 415472
rect 540720 411272 541520 411392
rect 0 403384 800 403504
rect 540720 399032 541520 399152
rect 0 391416 800 391536
rect 540720 386792 541520 386912
rect 0 379448 800 379568
rect 540720 374552 541520 374672
rect 0 367480 800 367600
rect 540720 362312 541520 362432
rect 0 355512 800 355632
rect 540720 350072 541520 350192
rect 0 343544 800 343664
rect 540720 337832 541520 337952
rect 0 331576 800 331696
rect 540720 325592 541520 325712
rect 0 319608 800 319728
rect 540720 313352 541520 313472
rect 0 307640 800 307760
rect 540720 301112 541520 301232
rect 0 295672 800 295792
rect 540720 288872 541520 288992
rect 0 283704 800 283824
rect 540720 276632 541520 276752
rect 0 271736 800 271856
rect 540720 264392 541520 264512
rect 0 259768 800 259888
rect 540720 252152 541520 252272
rect 0 247800 800 247920
rect 540720 239912 541520 240032
rect 0 235832 800 235952
rect 540720 227672 541520 227792
rect 0 223864 800 223984
rect 540720 215432 541520 215552
rect 0 211896 800 212016
rect 540720 203192 541520 203312
rect 0 199928 800 200048
rect 540720 190952 541520 191072
rect 0 187960 800 188080
rect 540720 178712 541520 178832
rect 0 175992 800 176112
rect 540720 166472 541520 166592
rect 0 164024 800 164144
rect 540720 154232 541520 154352
rect 0 152056 800 152176
rect 540720 141992 541520 142112
rect 0 140088 800 140208
rect 540720 129752 541520 129872
rect 0 128120 800 128240
rect 540720 117512 541520 117632
rect 0 116152 800 116272
rect 540720 105272 541520 105392
rect 0 104184 800 104304
rect 540720 93032 541520 93152
rect 0 92216 800 92336
rect 540720 80792 541520 80912
rect 0 80248 800 80368
rect 540720 68552 541520 68672
rect 0 68280 800 68400
rect 0 56312 800 56432
rect 540720 56312 541520 56432
rect 0 44344 800 44464
rect 540720 44072 541520 44192
rect 0 32376 800 32496
rect 540720 31832 541520 31952
rect 0 20408 800 20528
rect 540720 19592 541520 19712
rect 0 8440 800 8560
rect 540720 7352 541520 7472
<< obsm3 >>
rect 473 644032 541315 649025
rect 473 643752 540640 644032
rect 473 642944 541315 643752
rect 880 642664 541315 642944
rect 473 631792 541315 642664
rect 473 631512 540640 631792
rect 473 630976 541315 631512
rect 880 630696 541315 630976
rect 473 619552 541315 630696
rect 473 619272 540640 619552
rect 473 619008 541315 619272
rect 880 618728 541315 619008
rect 473 607312 541315 618728
rect 473 607040 540640 607312
rect 880 607032 540640 607040
rect 880 606760 541315 607032
rect 473 595072 541315 606760
rect 880 594792 540640 595072
rect 473 583104 541315 594792
rect 880 582832 541315 583104
rect 880 582824 540640 582832
rect 473 582552 540640 582824
rect 473 571136 541315 582552
rect 880 570856 541315 571136
rect 473 570592 541315 570856
rect 473 570312 540640 570592
rect 473 559168 541315 570312
rect 880 558888 541315 559168
rect 473 558352 541315 558888
rect 473 558072 540640 558352
rect 473 547200 541315 558072
rect 880 546920 541315 547200
rect 473 546112 541315 546920
rect 473 545832 540640 546112
rect 473 535232 541315 545832
rect 880 534952 541315 535232
rect 473 533872 541315 534952
rect 473 533592 540640 533872
rect 473 523264 541315 533592
rect 880 522984 541315 523264
rect 473 521632 541315 522984
rect 473 521352 540640 521632
rect 473 511296 541315 521352
rect 880 511016 541315 511296
rect 473 509392 541315 511016
rect 473 509112 540640 509392
rect 473 499328 541315 509112
rect 880 499048 541315 499328
rect 473 497152 541315 499048
rect 473 496872 540640 497152
rect 473 487360 541315 496872
rect 880 487080 541315 487360
rect 473 484912 541315 487080
rect 473 484632 540640 484912
rect 473 475392 541315 484632
rect 880 475112 541315 475392
rect 473 472672 541315 475112
rect 473 472392 540640 472672
rect 473 463424 541315 472392
rect 880 463144 541315 463424
rect 473 460432 541315 463144
rect 473 460152 540640 460432
rect 473 451456 541315 460152
rect 880 451176 541315 451456
rect 473 448192 541315 451176
rect 473 447912 540640 448192
rect 473 439488 541315 447912
rect 880 439208 541315 439488
rect 473 435952 541315 439208
rect 473 435672 540640 435952
rect 473 427520 541315 435672
rect 880 427240 541315 427520
rect 473 423712 541315 427240
rect 473 423432 540640 423712
rect 473 415552 541315 423432
rect 880 415272 541315 415552
rect 473 411472 541315 415272
rect 473 411192 540640 411472
rect 473 403584 541315 411192
rect 880 403304 541315 403584
rect 473 399232 541315 403304
rect 473 398952 540640 399232
rect 473 391616 541315 398952
rect 880 391336 541315 391616
rect 473 386992 541315 391336
rect 473 386712 540640 386992
rect 473 379648 541315 386712
rect 880 379368 541315 379648
rect 473 374752 541315 379368
rect 473 374472 540640 374752
rect 473 367680 541315 374472
rect 880 367400 541315 367680
rect 473 362512 541315 367400
rect 473 362232 540640 362512
rect 473 355712 541315 362232
rect 880 355432 541315 355712
rect 473 350272 541315 355432
rect 473 349992 540640 350272
rect 473 343744 541315 349992
rect 880 343464 541315 343744
rect 473 338032 541315 343464
rect 473 337752 540640 338032
rect 473 331776 541315 337752
rect 880 331496 541315 331776
rect 473 325792 541315 331496
rect 473 325512 540640 325792
rect 473 319808 541315 325512
rect 880 319528 541315 319808
rect 473 313552 541315 319528
rect 473 313272 540640 313552
rect 473 307840 541315 313272
rect 880 307560 541315 307840
rect 473 301312 541315 307560
rect 473 301032 540640 301312
rect 473 295872 541315 301032
rect 880 295592 541315 295872
rect 473 289072 541315 295592
rect 473 288792 540640 289072
rect 473 283904 541315 288792
rect 880 283624 541315 283904
rect 473 276832 541315 283624
rect 473 276552 540640 276832
rect 473 271936 541315 276552
rect 880 271656 541315 271936
rect 473 264592 541315 271656
rect 473 264312 540640 264592
rect 473 259968 541315 264312
rect 880 259688 541315 259968
rect 473 252352 541315 259688
rect 473 252072 540640 252352
rect 473 248000 541315 252072
rect 880 247720 541315 248000
rect 473 240112 541315 247720
rect 473 239832 540640 240112
rect 473 236032 541315 239832
rect 880 235752 541315 236032
rect 473 227872 541315 235752
rect 473 227592 540640 227872
rect 473 224064 541315 227592
rect 880 223784 541315 224064
rect 473 215632 541315 223784
rect 473 215352 540640 215632
rect 473 212096 541315 215352
rect 880 211816 541315 212096
rect 473 203392 541315 211816
rect 473 203112 540640 203392
rect 473 200128 541315 203112
rect 880 199848 541315 200128
rect 473 191152 541315 199848
rect 473 190872 540640 191152
rect 473 188160 541315 190872
rect 880 187880 541315 188160
rect 473 178912 541315 187880
rect 473 178632 540640 178912
rect 473 176192 541315 178632
rect 880 175912 541315 176192
rect 473 166672 541315 175912
rect 473 166392 540640 166672
rect 473 164224 541315 166392
rect 880 163944 541315 164224
rect 473 154432 541315 163944
rect 473 154152 540640 154432
rect 473 152256 541315 154152
rect 880 151976 541315 152256
rect 473 142192 541315 151976
rect 473 141912 540640 142192
rect 473 140288 541315 141912
rect 880 140008 541315 140288
rect 473 129952 541315 140008
rect 473 129672 540640 129952
rect 473 128320 541315 129672
rect 880 128040 541315 128320
rect 473 117712 541315 128040
rect 473 117432 540640 117712
rect 473 116352 541315 117432
rect 880 116072 541315 116352
rect 473 105472 541315 116072
rect 473 105192 540640 105472
rect 473 104384 541315 105192
rect 880 104104 541315 104384
rect 473 93232 541315 104104
rect 473 92952 540640 93232
rect 473 92416 541315 92952
rect 880 92136 541315 92416
rect 473 80992 541315 92136
rect 473 80712 540640 80992
rect 473 80448 541315 80712
rect 880 80168 541315 80448
rect 473 68752 541315 80168
rect 473 68480 540640 68752
rect 880 68472 540640 68480
rect 880 68200 541315 68472
rect 473 56512 541315 68200
rect 880 56232 540640 56512
rect 473 44544 541315 56232
rect 880 44272 541315 44544
rect 880 44264 540640 44272
rect 473 43992 540640 44264
rect 473 32576 541315 43992
rect 880 32296 541315 32576
rect 473 32032 541315 32296
rect 473 31752 540640 32032
rect 473 20608 541315 31752
rect 880 20328 541315 20608
rect 473 19792 541315 20328
rect 473 19512 540640 19792
rect 473 8640 541315 19512
rect 880 8360 541315 8640
rect 473 7552 541315 8360
rect 473 7272 540640 7552
rect 473 2143 541315 7272
<< metal4 >>
rect 4208 2128 4528 649040
rect 19568 2128 19888 649040
rect 34928 2128 35248 649040
rect 50288 2128 50608 649040
rect 65648 2128 65968 649040
rect 81008 2128 81328 649040
rect 96368 2128 96688 649040
rect 111728 2128 112048 649040
rect 127088 2128 127408 649040
rect 142448 2128 142768 649040
rect 157808 2128 158128 649040
rect 173168 2128 173488 649040
rect 188528 2128 188848 649040
rect 203888 2128 204208 649040
rect 219248 2128 219568 649040
rect 234608 2128 234928 649040
rect 249968 2128 250288 649040
rect 265328 2128 265648 649040
rect 280688 2128 281008 649040
rect 296048 2128 296368 649040
rect 311408 2128 311728 649040
rect 326768 2128 327088 649040
rect 342128 2128 342448 649040
rect 357488 2128 357808 649040
rect 372848 2128 373168 649040
rect 388208 2128 388528 649040
rect 403568 2128 403888 649040
rect 418928 2128 419248 649040
rect 434288 2128 434608 649040
rect 449648 2128 449968 649040
rect 465008 2128 465328 649040
rect 480368 2128 480688 649040
rect 495728 2128 496048 649040
rect 511088 2128 511408 649040
rect 526448 2128 526768 649040
<< obsm4 >>
rect 611 3163 4128 646101
rect 4608 3163 19488 646101
rect 19968 3163 34848 646101
rect 35328 3163 50208 646101
rect 50688 3163 65568 646101
rect 66048 3163 80928 646101
rect 81408 3163 96288 646101
rect 96768 3163 111648 646101
rect 112128 3163 127008 646101
rect 127488 3163 142368 646101
rect 142848 3163 157728 646101
rect 158208 3163 173088 646101
rect 173568 3163 188448 646101
rect 188928 3163 203808 646101
rect 204288 3163 219168 646101
rect 219648 3163 234528 646101
rect 235008 3163 249888 646101
rect 250368 3163 265248 646101
rect 265728 3163 280608 646101
rect 281088 3163 295968 646101
rect 296448 3163 311328 646101
rect 311808 3163 326688 646101
rect 327168 3163 342048 646101
rect 342528 3163 357408 646101
rect 357888 3163 372768 646101
rect 373248 3163 388128 646101
rect 388608 3163 403488 646101
rect 403968 3163 418848 646101
rect 419328 3163 434208 646101
rect 434688 3163 449568 646101
rect 450048 3163 464928 646101
rect 465408 3163 480288 646101
rect 480768 3163 495648 646101
rect 496128 3163 511008 646101
rect 511488 3163 526368 646101
rect 526848 3163 539797 646101
<< labels >>
rlabel metal3 s 540720 264392 541520 264512 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 413190 650726 413246 651526 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 353206 650726 353262 651526 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 293222 650726 293278 651526 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 233238 650726 233294 651526 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 173254 650726 173310 651526 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 113270 650726 113326 651526 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 53286 650726 53342 651526 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 642744 800 642864 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 594872 800 594992 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 547000 800 547120 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 540720 313352 541520 313472 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 499128 800 499248 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 451256 800 451376 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 403384 800 403504 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 0 355512 800 355632 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 307640 800 307760 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 259768 800 259888 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 211896 800 212016 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 164024 800 164144 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 0 116152 800 116272 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 540720 362312 541520 362432 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 540720 411272 541520 411392 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 540720 460232 541520 460352 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 540720 509192 541520 509312 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 540720 558152 541520 558272 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 540720 607112 541520 607232 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 533158 650726 533214 651526 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 473174 650726 473230 651526 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 540720 7352 541520 7472 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 540720 423512 541520 423632 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 540720 472472 541520 472592 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 540720 521432 541520 521552 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 540720 570392 541520 570512 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 540720 619352 541520 619472 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 518162 650726 518218 651526 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 458178 650726 458234 651526 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 398194 650726 398250 651526 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 338210 650726 338266 651526 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 278226 650726 278282 651526 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 540720 44072 541520 44192 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 218242 650726 218298 651526 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 158258 650726 158314 651526 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 98274 650726 98330 651526 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 38290 650726 38346 651526 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 630776 800 630896 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 0 582904 800 583024 6 io_in[25]
port 47 nsew signal input
rlabel metal3 s 0 535032 800 535152 6 io_in[26]
port 48 nsew signal input
rlabel metal3 s 0 487160 800 487280 6 io_in[27]
port 49 nsew signal input
rlabel metal3 s 0 439288 800 439408 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 391416 800 391536 6 io_in[29]
port 51 nsew signal input
rlabel metal3 s 540720 80792 541520 80912 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 0 343544 800 343664 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 0 295672 800 295792 6 io_in[31]
port 54 nsew signal input
rlabel metal3 s 0 247800 800 247920 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 199928 800 200048 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 0 152056 800 152176 6 io_in[34]
port 57 nsew signal input
rlabel metal3 s 0 104184 800 104304 6 io_in[35]
port 58 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 io_in[36]
port 59 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 io_in[37]
port 60 nsew signal input
rlabel metal3 s 540720 117512 541520 117632 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 540720 154232 541520 154352 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 540720 190952 541520 191072 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 540720 227672 541520 227792 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 540720 276632 541520 276752 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 540720 325592 541520 325712 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 540720 374552 541520 374672 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 540720 31832 541520 31952 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 540720 447992 541520 448112 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 540720 496952 541520 497072 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 540720 545912 541520 546032 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 540720 594872 541520 594992 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 540720 643832 541520 643952 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 488170 650726 488226 651526 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 428186 650726 428242 651526 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 368202 650726 368258 651526 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 308218 650726 308274 651526 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 248234 650726 248290 651526 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 540720 68552 541520 68672 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 188250 650726 188306 651526 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 128266 650726 128322 651526 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 68282 650726 68338 651526 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8298 650726 8354 651526 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 0 606840 800 606960 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 558968 800 559088 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 511096 800 511216 6 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s 0 463224 800 463344 6 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s 0 415352 800 415472 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 367480 800 367600 6 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 540720 105272 541520 105392 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 319608 800 319728 6 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s 0 271736 800 271856 6 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s 0 223864 800 223984 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 0 175992 800 176112 6 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s 0 128120 800 128240 6 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 540720 141992 541520 142112 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 540720 178712 541520 178832 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 540720 215432 541520 215552 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 540720 252152 541520 252272 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 540720 301112 541520 301232 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 540720 350072 541520 350192 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 540720 399032 541520 399152 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 540720 19592 541520 19712 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 540720 435752 541520 435872 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 540720 484712 541520 484832 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 540720 533672 541520 533792 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 540720 582632 541520 582752 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 540720 631592 541520 631712 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 503166 650726 503222 651526 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 443182 650726 443238 651526 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 383198 650726 383254 651526 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 323214 650726 323270 651526 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 263230 650726 263286 651526 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 540720 56312 541520 56432 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 203246 650726 203302 651526 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 143262 650726 143318 651526 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 83278 650726 83334 651526 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 23294 650726 23350 651526 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 0 618808 800 618928 6 io_out[24]
port 122 nsew signal output
rlabel metal3 s 0 570936 800 571056 6 io_out[25]
port 123 nsew signal output
rlabel metal3 s 0 523064 800 523184 6 io_out[26]
port 124 nsew signal output
rlabel metal3 s 0 475192 800 475312 6 io_out[27]
port 125 nsew signal output
rlabel metal3 s 0 427320 800 427440 6 io_out[28]
port 126 nsew signal output
rlabel metal3 s 0 379448 800 379568 6 io_out[29]
port 127 nsew signal output
rlabel metal3 s 540720 93032 541520 93152 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s 0 331576 800 331696 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 0 283704 800 283824 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 235832 800 235952 6 io_out[32]
port 131 nsew signal output
rlabel metal3 s 0 187960 800 188080 6 io_out[33]
port 132 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 io_out[35]
port 134 nsew signal output
rlabel metal3 s 0 56312 800 56432 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 io_out[37]
port 136 nsew signal output
rlabel metal3 s 540720 129752 541520 129872 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 540720 166472 541520 166592 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 540720 203192 541520 203312 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 540720 239912 541520 240032 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 540720 288872 541520 288992 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 540720 337832 541520 337952 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 540720 386792 541520 386912 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 128542 0 128598 800 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 432142 0 432198 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 435178 0 435234 800 6 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 438214 0 438270 800 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 441250 0 441306 800 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 444286 0 444342 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 447322 0 447378 800 6 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 450358 0 450414 800 6 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 453394 0 453450 800 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 456430 0 456486 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 459466 0 459522 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 462502 0 462558 800 6 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 465538 0 465594 800 6 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 468574 0 468630 800 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 471610 0 471666 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 474646 0 474702 800 6 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 477682 0 477738 800 6 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 480718 0 480774 800 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 483754 0 483810 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 486790 0 486846 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 489826 0 489882 800 6 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 161938 0 161994 800 6 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 492862 0 492918 800 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 495898 0 495954 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 498934 0 498990 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 501970 0 502026 800 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 505006 0 505062 800 6 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 508042 0 508098 800 6 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 511078 0 511134 800 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 514114 0 514170 800 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 177118 0 177174 800 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 180154 0 180210 800 6 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 183190 0 183246 800 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 186226 0 186282 800 6 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 189262 0 189318 800 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 192298 0 192354 800 6 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 195334 0 195390 800 6 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 198370 0 198426 800 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 201406 0 201462 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 204442 0 204498 800 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 207478 0 207534 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 210514 0 210570 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 213550 0 213606 800 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 216586 0 216642 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 219622 0 219678 800 6 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 222658 0 222714 800 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 228730 0 228786 800 6 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 231766 0 231822 800 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 234802 0 234858 800 6 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 237838 0 237894 800 6 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 240874 0 240930 800 6 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 243910 0 243966 800 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 246946 0 247002 800 6 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 249982 0 250038 800 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 253018 0 253074 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 256054 0 256110 800 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 259090 0 259146 800 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 262126 0 262182 800 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 265162 0 265218 800 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 268198 0 268254 800 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 271234 0 271290 800 6 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 274270 0 274326 800 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 277306 0 277362 800 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 280342 0 280398 800 6 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 283378 0 283434 800 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 286414 0 286470 800 6 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 289450 0 289506 800 6 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 292486 0 292542 800 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 295522 0 295578 800 6 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 298558 0 298614 800 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 301594 0 301650 800 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 304630 0 304686 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 307666 0 307722 800 6 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 310702 0 310758 800 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 313738 0 313794 800 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 316774 0 316830 800 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 319810 0 319866 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 322846 0 322902 800 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 325882 0 325938 800 6 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 328918 0 328974 800 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 331954 0 332010 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 334990 0 335046 800 6 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 338026 0 338082 800 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 341062 0 341118 800 6 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 344098 0 344154 800 6 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 347134 0 347190 800 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 350170 0 350226 800 6 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 353206 0 353262 800 6 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 356242 0 356298 800 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 359278 0 359334 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 362314 0 362370 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 365350 0 365406 800 6 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 368386 0 368442 800 6 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 371422 0 371478 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 374458 0 374514 800 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 377494 0 377550 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 380530 0 380586 800 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 383566 0 383622 800 6 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 386602 0 386658 800 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 389638 0 389694 800 6 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 392674 0 392730 800 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 395710 0 395766 800 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 398746 0 398802 800 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 401782 0 401838 800 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 404818 0 404874 800 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 407854 0 407910 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 410890 0 410946 800 6 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 413926 0 413982 800 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 416962 0 417018 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 419998 0 420054 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 423034 0 423090 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 426070 0 426126 800 6 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 429106 0 429162 800 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 433154 0 433210 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 436190 0 436246 800 6 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 439226 0 439282 800 6 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 442262 0 442318 800 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 445298 0 445354 800 6 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 448334 0 448390 800 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 451370 0 451426 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 454406 0 454462 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 457442 0 457498 800 6 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 460478 0 460534 800 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 159914 0 159970 800 6 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 463514 0 463570 800 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 466550 0 466606 800 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 469586 0 469642 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 472622 0 472678 800 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 475658 0 475714 800 6 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 478694 0 478750 800 6 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 481730 0 481786 800 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 484766 0 484822 800 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 487802 0 487858 800 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 490838 0 490894 800 6 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 493874 0 493930 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 496910 0 496966 800 6 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 499946 0 500002 800 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 502982 0 503038 800 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 506018 0 506074 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 509054 0 509110 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 512090 0 512146 800 6 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 515126 0 515182 800 6 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 165986 0 166042 800 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 169022 0 169078 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 172058 0 172114 800 6 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 175094 0 175150 800 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 178130 0 178186 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 181166 0 181222 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 184202 0 184258 800 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 187238 0 187294 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 132590 0 132646 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 190274 0 190330 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 193310 0 193366 800 6 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 196346 0 196402 800 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 199382 0 199438 800 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 202418 0 202474 800 6 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 205454 0 205510 800 6 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 208490 0 208546 800 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 211526 0 211582 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 214562 0 214618 800 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 217598 0 217654 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 135626 0 135682 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 220634 0 220690 800 6 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 223670 0 223726 800 6 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 226706 0 226762 800 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 229742 0 229798 800 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 232778 0 232834 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 235814 0 235870 800 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 238850 0 238906 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 241886 0 241942 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 244922 0 244978 800 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 247958 0 248014 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 138662 0 138718 800 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 250994 0 251050 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 254030 0 254086 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 257066 0 257122 800 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 260102 0 260158 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 263138 0 263194 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 266174 0 266230 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 269210 0 269266 800 6 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 272246 0 272302 800 6 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 275282 0 275338 800 6 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 278318 0 278374 800 6 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 281354 0 281410 800 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 284390 0 284446 800 6 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 287426 0 287482 800 6 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 290462 0 290518 800 6 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 293498 0 293554 800 6 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 296534 0 296590 800 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 299570 0 299626 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 302606 0 302662 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 305642 0 305698 800 6 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 308678 0 308734 800 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144734 0 144790 800 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 311714 0 311770 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 314750 0 314806 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 317786 0 317842 800 6 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 320822 0 320878 800 6 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 323858 0 323914 800 6 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 326894 0 326950 800 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 329930 0 329986 800 6 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 332966 0 333022 800 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 336002 0 336058 800 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 339038 0 339094 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 342074 0 342130 800 6 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 345110 0 345166 800 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 348146 0 348202 800 6 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 351182 0 351238 800 6 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 354218 0 354274 800 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 357254 0 357310 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 360290 0 360346 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 363326 0 363382 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 366362 0 366418 800 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 369398 0 369454 800 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 150806 0 150862 800 6 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 372434 0 372490 800 6 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 375470 0 375526 800 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 378506 0 378562 800 6 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 381542 0 381598 800 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 384578 0 384634 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 387614 0 387670 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 390650 0 390706 800 6 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 393686 0 393742 800 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 396722 0 396778 800 6 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 399758 0 399814 800 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 153842 0 153898 800 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 402794 0 402850 800 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 405830 0 405886 800 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 408866 0 408922 800 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 411902 0 411958 800 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 414938 0 414994 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 417974 0 418030 800 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 421010 0 421066 800 6 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 424046 0 424102 800 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 427082 0 427138 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 430118 0 430174 800 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 156878 0 156934 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 130566 0 130622 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 434166 0 434222 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 437202 0 437258 800 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 440238 0 440294 800 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 443274 0 443330 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 446310 0 446366 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 449346 0 449402 800 6 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 452382 0 452438 800 6 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 455418 0 455474 800 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 458454 0 458510 800 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 461490 0 461546 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 464526 0 464582 800 6 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 467562 0 467618 800 6 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 470598 0 470654 800 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 473634 0 473690 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 476670 0 476726 800 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 479706 0 479762 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 482742 0 482798 800 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 485778 0 485834 800 6 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 488814 0 488870 800 6 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 491850 0 491906 800 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 494886 0 494942 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 497922 0 497978 800 6 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 500958 0 501014 800 6 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 503994 0 504050 800 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 507030 0 507086 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 510066 0 510122 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 513102 0 513158 800 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 516138 0 516194 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 173070 0 173126 800 6 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 179142 0 179198 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 182178 0 182234 800 6 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 188250 0 188306 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 191286 0 191342 800 6 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 194322 0 194378 800 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 200394 0 200450 800 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 203430 0 203486 800 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 206466 0 206522 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 209502 0 209558 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 212538 0 212594 800 6 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 215574 0 215630 800 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 218610 0 218666 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 221646 0 221702 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 224682 0 224738 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 227718 0 227774 800 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 230754 0 230810 800 6 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 236826 0 236882 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 239862 0 239918 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 242898 0 242954 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 245934 0 245990 800 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 248970 0 249026 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 252006 0 252062 800 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 255042 0 255098 800 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 258078 0 258134 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 261114 0 261170 800 6 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 264150 0 264206 800 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 267186 0 267242 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 270222 0 270278 800 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 273258 0 273314 800 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 276294 0 276350 800 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 279330 0 279386 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 282366 0 282422 800 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 285402 0 285458 800 6 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 288438 0 288494 800 6 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 291474 0 291530 800 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 294510 0 294566 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 297546 0 297602 800 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 300582 0 300638 800 6 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 303618 0 303674 800 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 306654 0 306710 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 309690 0 309746 800 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 312726 0 312782 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 315762 0 315818 800 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 318798 0 318854 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 321834 0 321890 800 6 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 324870 0 324926 800 6 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 327906 0 327962 800 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 330942 0 330998 800 6 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 333978 0 334034 800 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 337014 0 337070 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 340050 0 340106 800 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 343086 0 343142 800 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 346122 0 346178 800 6 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 349158 0 349214 800 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 352194 0 352250 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 355230 0 355286 800 6 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 358266 0 358322 800 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 361302 0 361358 800 6 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 364338 0 364394 800 6 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 367374 0 367430 800 6 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 370410 0 370466 800 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 151818 0 151874 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 373446 0 373502 800 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 376482 0 376538 800 6 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 379518 0 379574 800 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 382554 0 382610 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 385590 0 385646 800 6 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 388626 0 388682 800 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 391662 0 391718 800 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 394698 0 394754 800 6 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 397734 0 397790 800 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 400770 0 400826 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 403806 0 403862 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 406842 0 406898 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 409878 0 409934 800 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 412914 0 412970 800 6 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 415950 0 416006 800 6 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 418986 0 419042 800 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 422022 0 422078 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 425058 0 425114 800 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 428094 0 428150 800 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 431130 0 431186 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 517150 0 517206 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 518162 0 518218 800 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 519174 0 519230 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 520186 0 520242 800 6 user_irq[2]
port 531 nsew signal output
rlabel metal4 s 4208 2128 4528 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 649040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 649040 6 vssd1
port 533 nsew ground bidirectional
rlabel metal2 s 21270 0 21326 800 6 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 91098 0 91154 800 6 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 94134 0 94190 800 6 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 103242 0 103298 800 6 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 109314 0 109370 800 6 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 121458 0 121514 800 6 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 541520 651526
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 729940544
string GDS_FILE /mnt/r/work/Rift2Go_2310_Sky130_MPW7/openlane/user_proj_example/runs/22_11_23_20_49/results/signoff/rift2Wrap.magic.gds
string GDS_START 2009388
<< end >>

