magic
tech sky130A
magscale 1 2
timestamp 1669311247
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 349154 700476 349160 700528
rect 349212 700516 349218 700528
rect 364978 700516 364984 700528
rect 349212 700488 364984 700516
rect 349212 700476 349218 700488
rect 364978 700476 364984 700488
rect 365036 700476 365042 700528
rect 514754 700408 514760 700460
rect 514812 700448 514818 700460
rect 543458 700448 543464 700460
rect 514812 700420 543464 700448
rect 514812 700408 514818 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 364334 700340 364340 700392
rect 364392 700380 364398 700392
rect 381170 700380 381176 700392
rect 364392 700352 381176 700380
rect 364392 700340 364398 700352
rect 381170 700340 381176 700352
rect 381228 700340 381234 700392
rect 394694 700340 394700 700392
rect 394752 700380 394758 700392
rect 413646 700380 413652 700392
rect 394752 700352 413652 700380
rect 394752 700340 394758 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 425054 700340 425060 700392
rect 425112 700380 425118 700392
rect 446122 700380 446128 700392
rect 425112 700352 446128 700380
rect 425112 700340 425118 700352
rect 446122 700340 446128 700352
rect 446180 700340 446186 700392
rect 454034 700340 454040 700392
rect 454092 700380 454098 700392
rect 478506 700380 478512 700392
rect 454092 700352 478512 700380
rect 454092 700340 454098 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 484394 700340 484400 700392
rect 484452 700380 484458 700392
rect 510982 700380 510988 700392
rect 484452 700352 510988 700380
rect 484452 700340 484458 700352
rect 510982 700340 510988 700352
rect 511040 700340 511046 700392
rect 529934 700340 529940 700392
rect 529992 700380 529998 700392
rect 559650 700380 559656 700392
rect 529992 700352 559656 700380
rect 529992 700340 529998 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 244274 700272 244280 700324
rect 244332 700312 244338 700324
rect 251450 700312 251456 700324
rect 244332 700284 251456 700312
rect 244332 700272 244338 700284
rect 251450 700272 251456 700284
rect 251508 700272 251514 700324
rect 274634 700272 274640 700324
rect 274692 700312 274698 700324
rect 283834 700312 283840 700324
rect 274692 700284 283840 700312
rect 274692 700272 274698 700284
rect 283834 700272 283840 700284
rect 283892 700272 283898 700324
rect 289814 700272 289820 700324
rect 289872 700312 289878 700324
rect 300118 700312 300124 700324
rect 289872 700284 300124 700312
rect 289872 700272 289878 700284
rect 300118 700272 300124 700284
rect 300176 700272 300182 700324
rect 304994 700272 305000 700324
rect 305052 700312 305058 700324
rect 316310 700312 316316 700324
rect 305052 700284 316316 700312
rect 305052 700272 305058 700284
rect 316310 700272 316316 700284
rect 316368 700272 316374 700324
rect 320174 700272 320180 700324
rect 320232 700312 320238 700324
rect 332502 700312 332508 700324
rect 320232 700284 332508 700312
rect 320232 700272 320238 700284
rect 332502 700272 332508 700284
rect 332560 700272 332566 700324
rect 333974 700272 333980 700324
rect 334032 700312 334038 700324
rect 348786 700312 348792 700324
rect 334032 700284 348792 700312
rect 334032 700272 334038 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 379514 700272 379520 700324
rect 379572 700312 379578 700324
rect 397454 700312 397460 700324
rect 379572 700284 397460 700312
rect 379572 700272 379578 700284
rect 397454 700272 397460 700284
rect 397512 700272 397518 700324
rect 409874 700272 409880 700324
rect 409932 700312 409938 700324
rect 429838 700312 429844 700324
rect 409932 700284 429844 700312
rect 409932 700272 409938 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 438854 700272 438860 700324
rect 438912 700312 438918 700324
rect 462314 700312 462320 700324
rect 438912 700284 462320 700312
rect 438912 700272 438918 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 469214 700272 469220 700324
rect 469272 700312 469278 700324
rect 494790 700312 494796 700324
rect 469272 700284 494796 700312
rect 469272 700272 469278 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 499574 700272 499580 700324
rect 499632 700312 499638 700324
rect 527174 700312 527180 700324
rect 499632 700284 527180 700312
rect 499632 700272 499638 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 545114 700272 545120 700324
rect 545172 700312 545178 700324
rect 575842 700312 575848 700324
rect 545172 700284 575848 700312
rect 545172 700272 545178 700284
rect 575842 700272 575848 700284
rect 575900 700272 575906 700324
rect 154114 699660 154120 699712
rect 154172 699700 154178 699712
rect 154574 699700 154580 699712
rect 154172 699672 154580 699700
rect 154172 699660 154178 699672
rect 154574 699660 154580 699672
rect 154632 699660 154638 699712
rect 213914 699660 213920 699712
rect 213972 699700 213978 699712
rect 218974 699700 218980 699712
rect 213972 699672 218980 699700
rect 213972 699660 213978 699672
rect 218974 699660 218980 699672
rect 219032 699660 219038 699712
rect 229094 699660 229100 699712
rect 229152 699700 229158 699712
rect 235166 699700 235172 699712
rect 229152 699672 235172 699700
rect 229152 699660 229158 699672
rect 235166 699660 235172 699672
rect 235224 699660 235230 699712
rect 259454 699660 259460 699712
rect 259512 699700 259518 699712
rect 267642 699700 267648 699712
rect 259512 699672 267648 699700
rect 259512 699660 259518 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 555418 696940 555424 696992
rect 555476 696980 555482 696992
rect 580166 696980 580172 696992
rect 555476 696952 580172 696980
rect 555476 696940 555482 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 555510 683136 555516 683188
rect 555568 683176 555574 683188
rect 580166 683176 580172 683188
rect 555568 683148 580172 683176
rect 555568 683136 555574 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 555602 670692 555608 670744
rect 555660 670732 555666 670744
rect 580166 670732 580172 670744
rect 555660 670704 580172 670732
rect 555660 670692 555666 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 104894 666476 104900 666528
rect 104952 666516 104958 666528
rect 109954 666516 109960 666528
rect 104952 666488 109960 666516
rect 104952 666476 104958 666488
rect 109954 666476 109960 666488
rect 110012 666476 110018 666528
rect 136634 666476 136640 666528
rect 136692 666516 136698 666528
rect 139946 666516 139952 666528
rect 136692 666488 139952 666516
rect 136692 666476 136698 666488
rect 139946 666476 139952 666488
rect 140004 666476 140010 666528
rect 200574 666476 200580 666528
rect 200632 666516 200638 666528
rect 201494 666516 201500 666528
rect 200632 666488 201500 666516
rect 200632 666476 200638 666488
rect 201494 666476 201500 666488
rect 201552 666476 201558 666528
rect 6914 665796 6920 665848
rect 6972 665836 6978 665848
rect 19978 665836 19984 665848
rect 6972 665808 19984 665836
rect 6972 665796 6978 665808
rect 19978 665796 19984 665808
rect 20036 665796 20042 665848
rect 23474 665796 23480 665848
rect 23532 665836 23538 665848
rect 34974 665836 34980 665848
rect 23532 665808 34980 665836
rect 23532 665796 23538 665808
rect 34974 665796 34980 665808
rect 35032 665796 35038 665848
rect 40034 665796 40040 665848
rect 40092 665836 40098 665848
rect 49970 665836 49976 665848
rect 40092 665808 49976 665836
rect 40092 665796 40098 665808
rect 49970 665796 49976 665808
rect 50028 665796 50034 665848
rect 56594 665796 56600 665848
rect 56652 665836 56658 665848
rect 64966 665836 64972 665848
rect 56652 665808 64972 665836
rect 56652 665796 56658 665808
rect 64966 665796 64972 665808
rect 65024 665796 65030 665848
rect 71774 665796 71780 665848
rect 71832 665836 71838 665848
rect 80054 665836 80060 665848
rect 71832 665808 80060 665836
rect 71832 665796 71838 665808
rect 80054 665796 80060 665808
rect 80112 665796 80118 665848
rect 185578 665660 185584 665712
rect 185636 665700 185642 665712
rect 186314 665700 186320 665712
rect 185636 665672 186320 665700
rect 185636 665660 185642 665672
rect 186314 665660 186320 665672
rect 186372 665660 186378 665712
rect 88334 665184 88340 665236
rect 88392 665224 88398 665236
rect 95234 665224 95240 665236
rect 88392 665196 95240 665224
rect 88392 665184 88398 665196
rect 95234 665184 95240 665196
rect 95292 665184 95298 665236
rect 121454 665184 121460 665236
rect 121512 665224 121518 665236
rect 124950 665224 124956 665236
rect 121512 665196 124956 665224
rect 121512 665184 121518 665196
rect 124950 665184 124956 665196
rect 125008 665184 125014 665236
rect 3418 655460 3424 655512
rect 3476 655500 3482 655512
rect 9398 655500 9404 655512
rect 3476 655472 9404 655500
rect 3476 655460 3482 655472
rect 9398 655460 9404 655472
rect 9456 655460 9462 655512
rect 555694 643084 555700 643136
rect 555752 643124 555758 643136
rect 580166 643124 580172 643136
rect 555752 643096 580172 643124
rect 555752 643084 555758 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3510 643016 3516 643068
rect 3568 643056 3574 643068
rect 9398 643056 9404 643068
rect 3568 643028 9404 643056
rect 3568 643016 3574 643028
rect 9398 643016 9404 643028
rect 9456 643016 9462 643068
rect 3602 632000 3608 632052
rect 3660 632040 3666 632052
rect 9398 632040 9404 632052
rect 3660 632012 9404 632040
rect 3660 632000 3666 632012
rect 9398 632000 9404 632012
rect 9456 632000 9462 632052
rect 555418 630640 555424 630692
rect 555476 630680 555482 630692
rect 579982 630680 579988 630692
rect 555476 630652 579988 630680
rect 555476 630640 555482 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 3694 619556 3700 619608
rect 3752 619596 3758 619608
rect 9398 619596 9404 619608
rect 3752 619568 9404 619596
rect 3752 619556 3758 619568
rect 9398 619556 9404 619568
rect 9456 619556 9462 619608
rect 555142 619556 555148 619608
rect 555200 619596 555206 619608
rect 580258 619596 580264 619608
rect 555200 619568 580264 619596
rect 555200 619556 555206 619568
rect 580258 619556 580264 619568
rect 580316 619556 580322 619608
rect 555510 616836 555516 616888
rect 555568 616876 555574 616888
rect 580166 616876 580172 616888
rect 555568 616848 580172 616876
rect 555568 616836 555574 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3418 607112 3424 607164
rect 3476 607152 3482 607164
rect 9398 607152 9404 607164
rect 3476 607124 9404 607152
rect 3476 607112 3482 607124
rect 9398 607112 9404 607124
rect 9456 607112 9462 607164
rect 555602 603100 555608 603152
rect 555660 603140 555666 603152
rect 580166 603140 580172 603152
rect 555660 603112 580172 603140
rect 555660 603100 555666 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 3510 596096 3516 596148
rect 3568 596136 3574 596148
rect 9398 596136 9404 596148
rect 3568 596108 9404 596136
rect 3568 596096 3574 596108
rect 9398 596096 9404 596108
rect 9456 596096 9462 596148
rect 555418 590656 555424 590708
rect 555476 590696 555482 590708
rect 579798 590696 579804 590708
rect 555476 590668 579804 590696
rect 555476 590656 555482 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3602 583652 3608 583704
rect 3660 583692 3666 583704
rect 9398 583692 9404 583704
rect 3660 583664 9404 583692
rect 3660 583652 3666 583664
rect 9398 583652 9404 583664
rect 9456 583652 9462 583704
rect 555510 576852 555516 576904
rect 555568 576892 555574 576904
rect 580166 576892 580172 576904
rect 555568 576864 580172 576892
rect 555568 576852 555574 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3694 571276 3700 571328
rect 3752 571316 3758 571328
rect 8662 571316 8668 571328
rect 3752 571288 8668 571316
rect 3752 571276 3758 571288
rect 8662 571276 8668 571288
rect 8720 571276 8726 571328
rect 555602 563048 555608 563100
rect 555660 563088 555666 563100
rect 579798 563088 579804 563100
rect 555660 563060 579804 563088
rect 555660 563048 555666 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 559648 3424 559700
rect 3476 559688 3482 559700
rect 9398 559688 9404 559700
rect 3476 559660 9404 559688
rect 3476 559648 3482 559660
rect 9398 559648 9404 559660
rect 9456 559648 9462 559700
rect 555418 550604 555424 550656
rect 555476 550644 555482 550656
rect 580166 550644 580172 550656
rect 555476 550616 580172 550644
rect 555476 550604 555482 550616
rect 580166 550604 580172 550616
rect 580224 550604 580230 550656
rect 3510 547816 3516 547868
rect 3568 547856 3574 547868
rect 8662 547856 8668 547868
rect 3568 547828 8668 547856
rect 3568 547816 3574 547828
rect 8662 547816 8668 547828
rect 8720 547816 8726 547868
rect 555694 536800 555700 536852
rect 555752 536840 555758 536852
rect 580166 536840 580172 536852
rect 555752 536812 580172 536840
rect 555752 536800 555758 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3602 535372 3608 535424
rect 3660 535412 3666 535424
rect 9398 535412 9404 535424
rect 3660 535384 9404 535412
rect 3660 535372 3666 535384
rect 9398 535372 9404 535384
rect 9456 535372 9462 535424
rect 555510 524424 555516 524476
rect 555568 524464 555574 524476
rect 580166 524464 580172 524476
rect 555568 524436 580172 524464
rect 555568 524424 555574 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 524356 3424 524408
rect 3476 524396 3482 524408
rect 9030 524396 9036 524408
rect 3476 524368 9036 524396
rect 3476 524356 3482 524368
rect 9030 524356 9036 524368
rect 9088 524356 9094 524408
rect 3510 511232 3516 511284
rect 3568 511272 3574 511284
rect 9398 511272 9404 511284
rect 3568 511244 9404 511272
rect 3568 511232 3574 511244
rect 9398 511232 9404 511244
rect 9456 511232 9462 511284
rect 555418 510620 555424 510672
rect 555476 510660 555482 510672
rect 580166 510660 580172 510672
rect 555476 510632 580172 510660
rect 555476 510620 555482 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3602 499468 3608 499520
rect 3660 499508 3666 499520
rect 9398 499508 9404 499520
rect 3660 499480 9404 499508
rect 3660 499468 3666 499480
rect 9398 499468 9404 499480
rect 9456 499468 9462 499520
rect 555602 496816 555608 496868
rect 555660 496856 555666 496868
rect 580166 496856 580172 496868
rect 555660 496828 580172 496856
rect 555660 496816 555666 496828
rect 580166 496816 580172 496828
rect 580224 496816 580230 496868
rect 3418 488452 3424 488504
rect 3476 488492 3482 488504
rect 9030 488492 9036 488504
rect 3476 488464 9036 488492
rect 3476 488452 3482 488464
rect 9030 488452 9036 488464
rect 9088 488452 9094 488504
rect 555510 484372 555516 484424
rect 555568 484412 555574 484424
rect 580166 484412 580172 484424
rect 555568 484384 580172 484412
rect 555568 484372 555574 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3694 476008 3700 476060
rect 3752 476048 3758 476060
rect 8662 476048 8668 476060
rect 3752 476020 8668 476048
rect 3752 476008 3758 476020
rect 8662 476008 8668 476020
rect 8720 476008 8726 476060
rect 555418 470568 555424 470620
rect 555476 470608 555482 470620
rect 579982 470608 579988 470620
rect 555476 470580 579988 470608
rect 555476 470568 555482 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 463020 3516 463072
rect 3568 463060 3574 463072
rect 9398 463060 9404 463072
rect 3568 463032 9404 463060
rect 3568 463020 3574 463032
rect 9398 463020 9404 463032
rect 9456 463020 9462 463072
rect 555510 456764 555516 456816
rect 555568 456804 555574 456816
rect 580166 456804 580172 456816
rect 555568 456776 580172 456804
rect 555568 456764 555574 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3602 452548 3608 452600
rect 3660 452588 3666 452600
rect 9030 452588 9036 452600
rect 3660 452560 9036 452588
rect 3660 452548 3666 452560
rect 9030 452548 9036 452560
rect 9088 452548 9094 452600
rect 555418 444388 555424 444440
rect 555476 444428 555482 444440
rect 580166 444428 580172 444440
rect 555476 444400 580172 444428
rect 555476 444388 555482 444400
rect 580166 444388 580172 444400
rect 580224 444388 580230 444440
rect 3418 440172 3424 440224
rect 3476 440212 3482 440224
rect 9398 440212 9404 440224
rect 3476 440184 9404 440212
rect 3476 440172 3482 440184
rect 9398 440172 9404 440184
rect 9456 440172 9462 440224
rect 555510 430584 555516 430636
rect 555568 430624 555574 430636
rect 580166 430624 580172 430636
rect 555568 430596 580172 430624
rect 555568 430584 555574 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3510 427728 3516 427780
rect 3568 427768 3574 427780
rect 9398 427768 9404 427780
rect 3568 427740 9404 427768
rect 3568 427728 3574 427740
rect 9398 427728 9404 427740
rect 9456 427728 9462 427780
rect 555418 418140 555424 418192
rect 555476 418180 555482 418192
rect 580166 418180 580172 418192
rect 555476 418152 580172 418180
rect 555476 418140 555482 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3418 416712 3424 416764
rect 3476 416752 3482 416764
rect 9030 416752 9036 416764
rect 3476 416724 9036 416752
rect 3476 416712 3482 416724
rect 9030 416712 9036 416724
rect 9088 416712 9094 416764
rect 555510 404336 555516 404388
rect 555568 404376 555574 404388
rect 580166 404376 580172 404388
rect 555568 404348 580172 404376
rect 555568 404336 555574 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 404268 3516 404320
rect 3568 404308 3574 404320
rect 9398 404308 9404 404320
rect 3568 404280 9404 404308
rect 3568 404268 3574 404280
rect 9398 404268 9404 404280
rect 9456 404268 9462 404320
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 7558 397508 7564 397520
rect 3568 397480 7564 397508
rect 3568 397468 3574 397480
rect 7558 397468 7564 397480
rect 7616 397468 7622 397520
rect 3418 391892 3424 391944
rect 3476 391932 3482 391944
rect 9398 391932 9404 391944
rect 3476 391904 9404 391932
rect 3476 391892 3482 391904
rect 9398 391892 9404 391904
rect 9456 391892 9462 391944
rect 555418 390532 555424 390584
rect 555476 390572 555482 390584
rect 580166 390572 580172 390584
rect 555476 390544 580172 390572
rect 555476 390532 555482 390544
rect 580166 390532 580172 390544
rect 580224 390532 580230 390584
rect 3418 383664 3424 383716
rect 3476 383704 3482 383716
rect 9030 383704 9036 383716
rect 3476 383676 9036 383704
rect 3476 383664 3482 383676
rect 9030 383664 9036 383676
rect 9088 383664 9094 383716
rect 555510 378156 555516 378208
rect 555568 378196 555574 378208
rect 580166 378196 580172 378208
rect 555568 378168 580172 378196
rect 555568 378156 555574 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3418 371288 3424 371340
rect 3476 371328 3482 371340
rect 8938 371328 8944 371340
rect 3476 371300 8944 371328
rect 3476 371288 3482 371300
rect 8938 371288 8944 371300
rect 8996 371288 9002 371340
rect 555602 364352 555608 364404
rect 555660 364392 555666 364404
rect 580166 364392 580172 364404
rect 555660 364364 580172 364392
rect 555660 364352 555666 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 2958 357416 2964 357468
rect 3016 357456 3022 357468
rect 6178 357456 6184 357468
rect 3016 357428 6184 357456
rect 3016 357416 3022 357428
rect 6178 357416 6184 357428
rect 6236 357416 6242 357468
rect 555418 351908 555424 351960
rect 555476 351948 555482 351960
rect 580166 351948 580172 351960
rect 555476 351920 580172 351948
rect 555476 351908 555482 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3418 345312 3424 345364
rect 3476 345352 3482 345364
rect 8938 345352 8944 345364
rect 3476 345324 8944 345352
rect 3476 345312 3482 345324
rect 8938 345312 8944 345324
rect 8996 345312 9002 345364
rect 6178 343544 6184 343596
rect 6236 343584 6242 343596
rect 9398 343584 9404 343596
rect 6236 343556 9404 343584
rect 6236 343544 6242 343556
rect 9398 343544 9404 343556
rect 9456 343544 9462 343596
rect 555510 338104 555516 338156
rect 555568 338144 555574 338156
rect 580166 338144 580172 338156
rect 555568 338116 580172 338144
rect 555568 338104 555574 338116
rect 580166 338104 580172 338116
rect 580224 338104 580230 338156
rect 3418 332256 3424 332308
rect 3476 332296 3482 332308
rect 7558 332296 7564 332308
rect 3476 332268 7564 332296
rect 3476 332256 3482 332268
rect 7558 332256 7564 332268
rect 7616 332256 7622 332308
rect 555418 324300 555424 324352
rect 555476 324340 555482 324352
rect 580166 324340 580172 324352
rect 555476 324312 580172 324340
rect 555476 324300 555482 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3418 319064 3424 319116
rect 3476 319104 3482 319116
rect 7650 319104 7656 319116
rect 3476 319076 7656 319104
rect 3476 319064 3482 319076
rect 7650 319064 7656 319076
rect 7708 319064 7714 319116
rect 555510 311856 555516 311908
rect 555568 311896 555574 311908
rect 580166 311896 580172 311908
rect 555568 311868 580172 311896
rect 555568 311856 555574 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 2774 305804 2780 305856
rect 2832 305844 2838 305856
rect 6178 305844 6184 305856
rect 2832 305816 6184 305844
rect 2832 305804 2838 305816
rect 6178 305804 6184 305816
rect 6236 305804 6242 305856
rect 555418 298120 555424 298172
rect 555476 298160 555482 298172
rect 580166 298160 580172 298172
rect 555476 298132 580172 298160
rect 555476 298120 555482 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 6178 296624 6184 296676
rect 6236 296664 6242 296676
rect 9490 296664 9496 296676
rect 6236 296636 9496 296664
rect 6236 296624 6242 296636
rect 9490 296624 9496 296636
rect 9548 296624 9554 296676
rect 2958 292544 2964 292596
rect 3016 292584 3022 292596
rect 6178 292584 6184 292596
rect 3016 292556 6184 292584
rect 3016 292544 3022 292556
rect 6178 292544 6184 292556
rect 6236 292544 6242 292596
rect 555418 284316 555424 284368
rect 555476 284356 555482 284368
rect 580166 284356 580172 284368
rect 555476 284328 580172 284356
rect 555476 284316 555482 284328
rect 580166 284316 580172 284328
rect 580224 284316 580230 284368
rect 6178 284248 6184 284300
rect 6236 284288 6242 284300
rect 8662 284288 8668 284300
rect 6236 284260 8668 284288
rect 6236 284248 6242 284260
rect 8662 284248 8668 284260
rect 8720 284248 8726 284300
rect 3510 279556 3516 279608
rect 3568 279596 3574 279608
rect 8202 279596 8208 279608
rect 3568 279568 8208 279596
rect 3568 279556 3574 279568
rect 8202 279556 8208 279568
rect 8260 279556 8266 279608
rect 555418 271872 555424 271924
rect 555476 271912 555482 271924
rect 579798 271912 579804 271924
rect 555476 271884 579804 271912
rect 555476 271872 555482 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 9398 266404 9404 266416
rect 3108 266376 9404 266404
rect 3108 266364 3114 266376
rect 9398 266364 9404 266376
rect 9456 266364 9462 266416
rect 556062 258068 556068 258120
rect 556120 258108 556126 258120
rect 580166 258108 580172 258120
rect 556120 258080 580172 258108
rect 556120 258068 556126 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 3418 254056 3424 254108
rect 3476 254096 3482 254108
rect 8938 254096 8944 254108
rect 3476 254068 8944 254096
rect 3476 254056 3482 254068
rect 8938 254056 8944 254068
rect 8996 254056 9002 254108
rect 555418 244264 555424 244316
rect 555476 244304 555482 244316
rect 579798 244304 579804 244316
rect 555476 244276 579804 244304
rect 555476 244264 555482 244276
rect 579798 244264 579804 244276
rect 579856 244264 579862 244316
rect 3694 235900 3700 235952
rect 3752 235940 3758 235952
rect 9398 235940 9404 235952
rect 3752 235912 9404 235940
rect 3752 235900 3758 235912
rect 9398 235900 9404 235912
rect 9456 235900 9462 235952
rect 555418 231820 555424 231872
rect 555476 231860 555482 231872
rect 580166 231860 580172 231872
rect 555476 231832 580172 231860
rect 555476 231820 555482 231832
rect 580166 231820 580172 231832
rect 580224 231820 580230 231872
rect 4154 224884 4160 224936
rect 4212 224924 4218 224936
rect 8846 224924 8852 224936
rect 4212 224896 8852 224924
rect 4212 224884 4218 224896
rect 8846 224884 8852 224896
rect 8904 224884 8910 224936
rect 555418 218016 555424 218068
rect 555476 218056 555482 218068
rect 580166 218056 580172 218068
rect 555476 218028 580172 218056
rect 555476 218016 555482 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 3142 213936 3148 213988
rect 3200 213976 3206 213988
rect 9214 213976 9220 213988
rect 3200 213948 9220 213976
rect 3200 213936 3206 213948
rect 9214 213936 9220 213948
rect 9272 213936 9278 213988
rect 555418 205640 555424 205692
rect 555476 205680 555482 205692
rect 580166 205680 580172 205692
rect 555476 205652 580172 205680
rect 555476 205640 555482 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 3418 201832 3424 201884
rect 3476 201872 3482 201884
rect 8294 201872 8300 201884
rect 3476 201844 8300 201872
rect 3476 201832 3482 201844
rect 8294 201832 8300 201844
rect 8352 201832 8358 201884
rect 580166 191876 580172 191888
rect 576826 191848 580172 191876
rect 555418 191768 555424 191820
rect 555476 191808 555482 191820
rect 576826 191808 576854 191848
rect 580166 191836 580172 191848
rect 580224 191836 580230 191888
rect 555476 191780 576854 191808
rect 555476 191768 555482 191780
rect 3418 188232 3424 188284
rect 3476 188272 3482 188284
rect 9398 188272 9404 188284
rect 3476 188244 9404 188272
rect 3476 188232 3482 188244
rect 9398 188232 9404 188244
rect 9456 188232 9462 188284
rect 555418 178644 555424 178696
rect 555476 178684 555482 178696
rect 580166 178684 580172 178696
rect 555476 178656 580172 178684
rect 555476 178644 555482 178656
rect 580166 178644 580172 178656
rect 580224 178644 580230 178696
rect 3326 175584 3332 175636
rect 3384 175624 3390 175636
rect 9398 175624 9404 175636
rect 3384 175596 9404 175624
rect 3384 175584 3390 175596
rect 9398 175584 9404 175596
rect 9456 175584 9462 175636
rect 555878 166268 555884 166320
rect 555936 166308 555942 166320
rect 580166 166308 580172 166320
rect 555936 166280 580172 166308
rect 555936 166268 555942 166280
rect 580166 166268 580172 166280
rect 580224 166268 580230 166320
rect 3418 162868 3424 162920
rect 3476 162908 3482 162920
rect 9398 162908 9404 162920
rect 3476 162880 9404 162908
rect 3476 162868 3482 162880
rect 9398 162868 9404 162880
rect 9456 162868 9462 162920
rect 555418 153212 555424 153264
rect 555476 153252 555482 153264
rect 579522 153252 579528 153264
rect 555476 153224 579528 153252
rect 555476 153212 555482 153224
rect 579522 153212 579528 153224
rect 579580 153212 579586 153264
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 8202 150396 8208 150408
rect 3476 150368 8208 150396
rect 3476 150356 3482 150368
rect 8202 150356 8208 150368
rect 8260 150356 8266 150408
rect 555418 139340 555424 139392
rect 555476 139380 555482 139392
rect 580166 139380 580172 139392
rect 555476 139352 580172 139380
rect 555476 139340 555482 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3234 136960 3240 137012
rect 3292 137000 3298 137012
rect 8202 137000 8208 137012
rect 3292 136972 8208 137000
rect 3292 136960 3298 136972
rect 8202 136960 8208 136972
rect 8260 136960 8266 137012
rect 555418 126896 555424 126948
rect 555476 126936 555482 126948
rect 580166 126936 580172 126948
rect 555476 126908 580172 126936
rect 555476 126896 555482 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 3418 123836 3424 123888
rect 3476 123876 3482 123888
rect 8202 123876 8208 123888
rect 3476 123848 8208 123876
rect 3476 123836 3482 123848
rect 8202 123836 8208 123848
rect 8260 123836 8266 123888
rect 555418 113092 555424 113144
rect 555476 113132 555482 113144
rect 579798 113132 579804 113144
rect 555476 113104 579804 113132
rect 555476 113092 555482 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3418 110712 3424 110764
rect 3476 110752 3482 110764
rect 8938 110752 8944 110764
rect 3476 110724 8944 110752
rect 3476 110712 3482 110724
rect 8938 110712 8944 110724
rect 8996 110712 9002 110764
rect 4154 103504 4160 103556
rect 4212 103544 4218 103556
rect 9398 103544 9404 103556
rect 4212 103516 9404 103544
rect 4212 103504 4218 103516
rect 9398 103504 9404 103516
rect 9456 103504 9462 103556
rect 555694 100648 555700 100700
rect 555752 100688 555758 100700
rect 580166 100688 580172 100700
rect 555752 100660 580172 100688
rect 555752 100648 555758 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 4154 91060 4160 91112
rect 4212 91100 4218 91112
rect 9398 91100 9404 91112
rect 4212 91072 9404 91100
rect 4212 91060 4218 91072
rect 9398 91060 9404 91072
rect 9456 91060 9462 91112
rect 554774 86912 554780 86964
rect 554832 86952 554838 86964
rect 580166 86952 580172 86964
rect 554832 86924 580172 86952
rect 554832 86912 554838 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 555418 73108 555424 73160
rect 555476 73148 555482 73160
rect 580166 73148 580172 73160
rect 555476 73120 580172 73148
rect 555476 73108 555482 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3418 71612 3424 71664
rect 3476 71652 3482 71664
rect 8938 71652 8944 71664
rect 3476 71624 8944 71652
rect 3476 71612 3482 71624
rect 8938 71612 8944 71624
rect 8996 71612 9002 71664
rect 555418 60664 555424 60716
rect 555476 60704 555482 60716
rect 580166 60704 580172 60716
rect 555476 60676 580172 60704
rect 555476 60664 555482 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3142 59168 3148 59220
rect 3200 59208 3206 59220
rect 8938 59208 8944 59220
rect 3200 59180 8944 59208
rect 3200 59168 3206 59180
rect 8938 59168 8944 59180
rect 8996 59168 9002 59220
rect 4798 55224 4804 55276
rect 4856 55264 4862 55276
rect 9398 55264 9404 55276
rect 4856 55236 9404 55264
rect 4856 55224 4862 55236
rect 9398 55224 9404 55236
rect 9456 55224 9462 55276
rect 555418 46860 555424 46912
rect 555476 46900 555482 46912
rect 580166 46900 580172 46912
rect 555476 46872 580172 46900
rect 555476 46860 555482 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 2774 45500 2780 45552
rect 2832 45540 2838 45552
rect 4798 45540 4804 45552
rect 2832 45512 4804 45540
rect 2832 45500 2838 45512
rect 4798 45500 4804 45512
rect 4856 45500 4862 45552
rect 3418 44140 3424 44192
rect 3476 44180 3482 44192
rect 9398 44180 9404 44192
rect 3476 44152 9404 44180
rect 3476 44140 3482 44152
rect 9398 44140 9404 44152
rect 9456 44140 9462 44192
rect 555418 33056 555424 33108
rect 555476 33096 555482 33108
rect 580166 33096 580172 33108
rect 555476 33068 580172 33096
rect 555476 33056 555482 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3510 31764 3516 31816
rect 3568 31804 3574 31816
rect 9398 31804 9404 31816
rect 3568 31776 9404 31804
rect 3568 31764 3574 31776
rect 9398 31764 9404 31776
rect 9456 31764 9462 31816
rect 555510 20612 555516 20664
rect 555568 20652 555574 20664
rect 579982 20652 579988 20664
rect 555568 20624 579988 20652
rect 555568 20612 555574 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 6178 19320 6184 19372
rect 6236 19360 6242 19372
rect 9398 19360 9404 19372
rect 6236 19332 9404 19360
rect 6236 19320 6242 19332
rect 9398 19320 9404 19332
rect 9456 19320 9462 19372
rect 219434 9596 219440 9648
rect 219492 9636 219498 9648
rect 220170 9636 220176 9648
rect 219492 9608 220176 9636
rect 219492 9596 219498 9608
rect 220170 9596 220176 9608
rect 220228 9596 220234 9648
rect 322842 9596 322848 9648
rect 322900 9636 322906 9648
rect 335538 9636 335544 9648
rect 322900 9608 335544 9636
rect 322900 9596 322906 9608
rect 335538 9596 335544 9608
rect 335596 9596 335602 9648
rect 340230 9596 340236 9648
rect 340288 9636 340294 9648
rect 356330 9636 356336 9648
rect 340288 9608 356336 9636
rect 340288 9596 340294 9608
rect 356330 9596 356336 9608
rect 356388 9596 356394 9648
rect 492030 9596 492036 9648
rect 492088 9636 492094 9648
rect 498194 9636 498200 9648
rect 492088 9608 498200 9636
rect 492088 9596 492094 9608
rect 498194 9596 498200 9608
rect 498252 9596 498258 9648
rect 499574 9596 499580 9648
rect 499632 9636 499638 9648
rect 500494 9636 500500 9648
rect 499632 9608 500500 9636
rect 499632 9596 499638 9608
rect 500494 9596 500500 9608
rect 500552 9596 500558 9648
rect 143626 9528 143632 9580
rect 143684 9568 143690 9580
rect 150434 9568 150440 9580
rect 143684 9540 150440 9568
rect 143684 9528 143690 9540
rect 150434 9528 150440 9540
rect 150492 9528 150498 9580
rect 151906 9528 151912 9580
rect 151964 9568 151970 9580
rect 157426 9568 157432 9580
rect 151964 9540 157432 9568
rect 151964 9528 151970 9540
rect 157426 9528 157432 9540
rect 157484 9528 157490 9580
rect 165982 9528 165988 9580
rect 166040 9568 166046 9580
rect 168558 9568 168564 9580
rect 166040 9540 168564 9568
rect 166040 9528 166046 9540
rect 168558 9528 168564 9540
rect 168616 9528 168622 9580
rect 261294 9528 261300 9580
rect 261352 9568 261358 9580
rect 263502 9568 263508 9580
rect 261352 9540 263508 9568
rect 261352 9528 261358 9540
rect 263502 9528 263508 9540
rect 263560 9528 263566 9580
rect 307662 9528 307668 9580
rect 307720 9568 307726 9580
rect 307720 9540 309824 9568
rect 307720 9528 307726 9540
rect 33134 9460 33140 9512
rect 33192 9500 33198 9512
rect 33962 9500 33968 9512
rect 33192 9472 33968 9500
rect 33192 9460 33198 9472
rect 33962 9460 33968 9472
rect 34020 9460 34026 9512
rect 44174 9460 44180 9512
rect 44232 9500 44238 9512
rect 45094 9500 45100 9512
rect 44232 9472 45100 9500
rect 44232 9460 44238 9472
rect 45094 9460 45100 9472
rect 45152 9460 45158 9512
rect 55214 9460 55220 9512
rect 55272 9500 55278 9512
rect 56226 9500 56232 9512
rect 55272 9472 56232 9500
rect 55272 9460 55278 9472
rect 56226 9460 56232 9472
rect 56284 9460 56290 9512
rect 67634 9460 67640 9512
rect 67692 9500 67698 9512
rect 68370 9500 68376 9512
rect 67692 9472 68376 9500
rect 67692 9460 67698 9472
rect 68370 9460 68376 9472
rect 68428 9460 68434 9512
rect 70394 9460 70400 9512
rect 70452 9500 70458 9512
rect 71406 9500 71412 9512
rect 70452 9472 71412 9500
rect 70452 9460 70458 9472
rect 71406 9460 71412 9472
rect 71464 9460 71470 9512
rect 85574 9460 85580 9512
rect 85632 9500 85638 9512
rect 86586 9500 86592 9512
rect 85632 9472 86592 9500
rect 85632 9460 85638 9472
rect 86586 9460 86592 9472
rect 86644 9460 86650 9512
rect 89714 9460 89720 9512
rect 89772 9500 89778 9512
rect 90634 9500 90640 9512
rect 89772 9472 90640 9500
rect 89772 9460 89778 9472
rect 90634 9460 90640 9472
rect 90692 9460 90698 9512
rect 107654 9460 107660 9512
rect 107712 9500 107718 9512
rect 109862 9500 109868 9512
rect 107712 9472 109868 9500
rect 107712 9460 107718 9472
rect 109862 9460 109868 9472
rect 109920 9460 109926 9512
rect 110322 9460 110328 9512
rect 110380 9500 110386 9512
rect 110874 9500 110880 9512
rect 110380 9472 110880 9500
rect 110380 9460 110386 9472
rect 110874 9460 110880 9472
rect 110932 9460 110938 9512
rect 116946 9460 116952 9512
rect 117004 9500 117010 9512
rect 120074 9500 120080 9512
rect 117004 9472 120080 9500
rect 117004 9460 117010 9472
rect 120074 9460 120080 9472
rect 120132 9460 120138 9512
rect 121362 9460 121368 9512
rect 121420 9500 121426 9512
rect 122006 9500 122012 9512
rect 121420 9472 122012 9500
rect 121420 9460 121426 9472
rect 122006 9460 122012 9472
rect 122064 9460 122070 9512
rect 131022 9460 131028 9512
rect 131080 9500 131086 9512
rect 132126 9500 132132 9512
rect 131080 9472 132132 9500
rect 131080 9460 131086 9472
rect 132126 9460 132132 9472
rect 132184 9460 132190 9512
rect 133966 9460 133972 9512
rect 134024 9500 134030 9512
rect 141234 9500 141240 9512
rect 134024 9472 141240 9500
rect 134024 9460 134030 9472
rect 141234 9460 141240 9472
rect 141292 9460 141298 9512
rect 146202 9460 146208 9512
rect 146260 9500 146266 9512
rect 151354 9500 151360 9512
rect 146260 9472 151360 9500
rect 146260 9460 146266 9472
rect 151354 9460 151360 9472
rect 151412 9460 151418 9512
rect 157242 9460 157248 9512
rect 157300 9500 157306 9512
rect 160462 9500 160468 9512
rect 157300 9472 160468 9500
rect 157300 9460 157306 9472
rect 160462 9460 160468 9472
rect 160520 9460 160526 9512
rect 167270 9460 167276 9512
rect 167328 9500 167334 9512
rect 169754 9500 169760 9512
rect 167328 9472 169760 9500
rect 167328 9460 167334 9472
rect 169754 9460 169760 9472
rect 169812 9460 169818 9512
rect 171226 9460 171232 9512
rect 171284 9500 171290 9512
rect 173894 9500 173900 9512
rect 171284 9472 173900 9500
rect 171284 9460 171290 9472
rect 173894 9460 173900 9472
rect 173952 9460 173958 9512
rect 175274 9460 175280 9512
rect 175332 9500 175338 9512
rect 177666 9500 177672 9512
rect 175332 9472 177672 9500
rect 175332 9460 175338 9472
rect 177666 9460 177672 9472
rect 177724 9460 177730 9512
rect 200114 9460 200120 9512
rect 200172 9500 200178 9512
rect 200942 9500 200948 9512
rect 200172 9472 200948 9500
rect 200172 9460 200178 9472
rect 200942 9460 200948 9472
rect 201000 9460 201006 9512
rect 201494 9460 201500 9512
rect 201552 9500 201558 9512
rect 204990 9500 204996 9512
rect 201552 9472 204996 9500
rect 201552 9460 201558 9472
rect 204990 9460 204996 9472
rect 205048 9460 205054 9512
rect 206186 9460 206192 9512
rect 206244 9500 206250 9512
rect 209038 9500 209044 9512
rect 206244 9472 209044 9500
rect 206244 9460 206250 9472
rect 209038 9460 209044 9472
rect 209096 9460 209102 9512
rect 210970 9460 210976 9512
rect 211028 9500 211034 9512
rect 213086 9500 213092 9512
rect 211028 9472 213092 9500
rect 211028 9460 211034 9472
rect 213086 9460 213092 9472
rect 213144 9460 213150 9512
rect 213362 9460 213368 9512
rect 213420 9500 213426 9512
rect 215294 9500 215300 9512
rect 213420 9472 215300 9500
rect 213420 9460 213426 9472
rect 215294 9460 215300 9472
rect 215352 9460 215358 9512
rect 215662 9460 215668 9512
rect 215720 9500 215726 9512
rect 217134 9500 217140 9512
rect 215720 9472 217140 9500
rect 215720 9460 215726 9472
rect 217134 9460 217140 9472
rect 217192 9460 217198 9512
rect 231762 9460 231768 9512
rect 231820 9500 231826 9512
rect 232222 9500 232228 9512
rect 231820 9472 232228 9500
rect 231820 9460 231826 9472
rect 232222 9460 232228 9472
rect 232280 9460 232286 9512
rect 232958 9460 232964 9512
rect 233016 9500 233022 9512
rect 233418 9500 233424 9512
rect 233016 9472 233424 9500
rect 233016 9460 233022 9472
rect 233418 9460 233424 9472
rect 233476 9460 233482 9512
rect 233970 9460 233976 9512
rect 234028 9500 234034 9512
rect 234706 9500 234712 9512
rect 234028 9472 234712 9500
rect 234028 9460 234034 9472
rect 234706 9460 234712 9472
rect 234764 9460 234770 9512
rect 235902 9460 235908 9512
rect 235960 9500 235966 9512
rect 237006 9500 237012 9512
rect 235960 9472 237012 9500
rect 235960 9460 235966 9472
rect 237006 9460 237012 9472
rect 237064 9460 237070 9512
rect 245102 9460 245108 9512
rect 245160 9500 245166 9512
rect 245838 9500 245844 9512
rect 245160 9472 245844 9500
rect 245160 9460 245166 9472
rect 245838 9460 245844 9472
rect 245896 9460 245902 9512
rect 251082 9460 251088 9512
rect 251140 9500 251146 9512
rect 252278 9500 252284 9512
rect 251140 9472 252284 9500
rect 251140 9460 251146 9472
rect 252278 9460 252284 9472
rect 252336 9460 252342 9512
rect 253842 9460 253848 9512
rect 253900 9500 253906 9512
rect 255222 9500 255228 9512
rect 253900 9472 255228 9500
rect 253900 9460 253906 9472
rect 255222 9460 255228 9472
rect 255280 9460 255286 9512
rect 256234 9460 256240 9512
rect 256292 9500 256298 9512
rect 257890 9500 257896 9512
rect 256292 9472 257896 9500
rect 256292 9460 256298 9472
rect 257890 9460 257896 9472
rect 257948 9460 257954 9512
rect 262122 9460 262128 9512
rect 262180 9500 262186 9512
rect 263410 9500 263416 9512
rect 262180 9472 263416 9500
rect 262180 9460 262186 9472
rect 263410 9460 263416 9472
rect 263468 9460 263474 9512
rect 265342 9460 265348 9512
rect 265400 9500 265406 9512
rect 267642 9500 267648 9512
rect 265400 9472 267648 9500
rect 265400 9460 265406 9472
rect 267642 9460 267648 9472
rect 267700 9460 267706 9512
rect 273070 9460 273076 9512
rect 273128 9500 273134 9512
rect 274542 9500 274548 9512
rect 273128 9472 274548 9500
rect 273128 9460 273134 9472
rect 274542 9460 274548 9472
rect 274600 9460 274606 9512
rect 275462 9460 275468 9512
rect 275520 9500 275526 9512
rect 276750 9500 276756 9512
rect 275520 9472 276756 9500
rect 275520 9460 275526 9472
rect 276750 9460 276756 9472
rect 276808 9460 276814 9512
rect 280522 9460 280528 9512
rect 280580 9500 280586 9512
rect 282822 9500 282828 9512
rect 280580 9472 282828 9500
rect 280580 9460 280586 9472
rect 282822 9460 282828 9472
rect 282880 9460 282886 9512
rect 283558 9460 283564 9512
rect 283616 9500 283622 9512
rect 285490 9500 285496 9512
rect 283616 9472 285496 9500
rect 283616 9460 283622 9472
rect 285490 9460 285496 9472
rect 285548 9460 285554 9512
rect 287606 9460 287612 9512
rect 287664 9500 287670 9512
rect 288526 9500 288532 9512
rect 287664 9472 288532 9500
rect 287664 9460 287670 9472
rect 288526 9460 288532 9472
rect 288584 9460 288590 9512
rect 292482 9460 292488 9512
rect 292540 9500 292546 9512
rect 293862 9500 293868 9512
rect 292540 9472 293868 9500
rect 292540 9460 292546 9472
rect 293862 9460 293868 9472
rect 293920 9460 293926 9512
rect 301774 9460 301780 9512
rect 301832 9500 301838 9512
rect 303062 9500 303068 9512
rect 301832 9472 303068 9500
rect 301832 9460 301838 9472
rect 303062 9460 303068 9472
rect 303120 9460 303126 9512
rect 306834 9460 306840 9512
rect 306892 9500 306898 9512
rect 308030 9500 308036 9512
rect 306892 9472 308036 9500
rect 306892 9460 306898 9472
rect 308030 9460 308036 9472
rect 308088 9460 308094 9512
rect 309796 9500 309824 9540
rect 309870 9528 309876 9580
rect 309928 9568 309934 9580
rect 316034 9568 316040 9580
rect 309928 9540 316040 9568
rect 309928 9528 309934 9540
rect 316034 9528 316040 9540
rect 316092 9528 316098 9580
rect 319990 9528 319996 9580
rect 320048 9568 320054 9580
rect 320048 9540 326016 9568
rect 320048 9528 320054 9540
rect 320910 9500 320916 9512
rect 309796 9472 316034 9500
rect 63402 9392 63408 9444
rect 63460 9432 63466 9444
rect 64322 9432 64328 9444
rect 63460 9404 64328 9432
rect 63460 9392 63466 9404
rect 64322 9392 64328 9404
rect 64380 9392 64386 9444
rect 97902 9392 97908 9444
rect 97960 9432 97966 9444
rect 98730 9432 98736 9444
rect 97960 9404 98736 9432
rect 97960 9392 97966 9404
rect 98730 9392 98736 9404
rect 98788 9392 98794 9444
rect 140866 9392 140872 9444
rect 140924 9432 140930 9444
rect 147306 9432 147312 9444
rect 140924 9404 147312 9432
rect 140924 9392 140930 9404
rect 147306 9392 147312 9404
rect 147364 9392 147370 9444
rect 153194 9392 153200 9444
rect 153252 9432 153258 9444
rect 158714 9432 158720 9444
rect 153252 9404 158720 9432
rect 153252 9392 153258 9404
rect 158714 9392 158720 9404
rect 158772 9392 158778 9444
rect 165338 9392 165344 9444
rect 165396 9432 165402 9444
rect 167546 9432 167552 9444
rect 165396 9404 167552 9432
rect 165396 9392 165402 9404
rect 167546 9392 167552 9404
rect 167604 9392 167610 9444
rect 175182 9392 175188 9444
rect 175240 9432 175246 9444
rect 175642 9432 175648 9444
rect 175240 9404 175648 9432
rect 175240 9392 175246 9404
rect 175642 9392 175648 9404
rect 175700 9392 175706 9444
rect 221550 9392 221556 9444
rect 221608 9432 221614 9444
rect 222194 9432 222200 9444
rect 221608 9404 222200 9432
rect 221608 9392 221614 9404
rect 222194 9392 222200 9404
rect 222252 9392 222258 9444
rect 236914 9392 236920 9444
rect 236972 9432 236978 9444
rect 238110 9432 238116 9444
rect 236972 9404 238116 9432
rect 236972 9392 236978 9404
rect 238110 9392 238116 9404
rect 238168 9392 238174 9444
rect 246942 9392 246948 9444
rect 247000 9432 247006 9444
rect 247862 9432 247868 9444
rect 247000 9404 247868 9432
rect 247000 9392 247006 9404
rect 247862 9392 247868 9404
rect 247920 9392 247926 9444
rect 252186 9392 252192 9444
rect 252244 9432 252250 9444
rect 253474 9432 253480 9444
rect 252244 9404 253480 9432
rect 252244 9392 252250 9404
rect 253474 9392 253480 9404
rect 253532 9392 253538 9444
rect 263318 9392 263324 9444
rect 263376 9432 263382 9444
rect 264882 9432 264888 9444
rect 263376 9404 264888 9432
rect 263376 9392 263382 9404
rect 264882 9392 264888 9404
rect 264940 9392 264946 9444
rect 274450 9392 274456 9444
rect 274508 9432 274514 9444
rect 275830 9432 275836 9444
rect 274508 9404 275836 9432
rect 274508 9392 274514 9404
rect 275830 9392 275836 9404
rect 275888 9392 275894 9444
rect 285582 9392 285588 9444
rect 285640 9432 285646 9444
rect 286134 9432 286140 9444
rect 285640 9404 286140 9432
rect 285640 9392 285646 9404
rect 286134 9392 286140 9404
rect 286192 9392 286198 9444
rect 294690 9392 294696 9444
rect 294748 9432 294754 9444
rect 295886 9432 295892 9444
rect 294748 9404 295892 9432
rect 294748 9392 294754 9404
rect 295886 9392 295892 9404
rect 295944 9392 295950 9444
rect 300762 9392 300768 9444
rect 300820 9432 300826 9444
rect 302142 9432 302148 9444
rect 300820 9404 302148 9432
rect 300820 9392 300826 9404
rect 302142 9392 302148 9404
rect 302200 9392 302206 9444
rect 304810 9392 304816 9444
rect 304868 9432 304874 9444
rect 305914 9432 305920 9444
rect 304868 9404 305920 9432
rect 304868 9392 304874 9404
rect 305914 9392 305920 9404
rect 305972 9392 305978 9444
rect 316006 9432 316034 9472
rect 316420 9472 320916 9500
rect 316420 9432 316448 9472
rect 320910 9460 320916 9472
rect 320968 9460 320974 9512
rect 321002 9460 321008 9512
rect 321060 9500 321066 9512
rect 325878 9500 325884 9512
rect 321060 9472 325884 9500
rect 321060 9460 321066 9472
rect 325878 9460 325884 9472
rect 325936 9460 325942 9512
rect 325988 9500 326016 9540
rect 326062 9528 326068 9580
rect 326120 9568 326126 9580
rect 340414 9568 340420 9580
rect 326120 9540 340420 9568
rect 326120 9528 326126 9540
rect 340414 9528 340420 9540
rect 340472 9528 340478 9580
rect 341242 9528 341248 9580
rect 341300 9568 341306 9580
rect 359918 9568 359924 9580
rect 341300 9540 359924 9568
rect 341300 9528 341306 9540
rect 359918 9528 359924 9540
rect 359976 9528 359982 9580
rect 496722 9528 496728 9580
rect 496780 9568 496786 9580
rect 525426 9568 525432 9580
rect 496780 9540 525432 9568
rect 496780 9528 496786 9540
rect 525426 9528 525432 9540
rect 525484 9528 525490 9580
rect 327994 9500 328000 9512
rect 325988 9472 328000 9500
rect 327994 9460 328000 9472
rect 328052 9460 328058 9512
rect 328086 9460 328092 9512
rect 328144 9500 328150 9512
rect 334066 9500 334072 9512
rect 328144 9472 334072 9500
rect 328144 9460 328150 9472
rect 334066 9460 334072 9472
rect 334124 9460 334130 9512
rect 343266 9460 343272 9512
rect 343324 9500 343330 9512
rect 343726 9500 343732 9512
rect 343324 9472 343732 9500
rect 343324 9460 343330 9472
rect 343726 9460 343732 9472
rect 343784 9460 343790 9512
rect 344278 9460 344284 9512
rect 344336 9500 344342 9512
rect 361758 9500 361764 9512
rect 344336 9472 361764 9500
rect 344336 9460 344342 9472
rect 361758 9460 361764 9472
rect 361816 9460 361822 9512
rect 366542 9460 366548 9512
rect 366600 9500 366606 9512
rect 371878 9500 371884 9512
rect 366600 9472 371884 9500
rect 366600 9460 366606 9472
rect 371878 9460 371884 9472
rect 371936 9460 371942 9512
rect 378134 9460 378140 9512
rect 378192 9500 378198 9512
rect 379054 9500 379060 9512
rect 378192 9472 379060 9500
rect 378192 9460 378198 9472
rect 379054 9460 379060 9472
rect 379112 9460 379118 9512
rect 404998 9460 405004 9512
rect 405056 9500 405062 9512
rect 406378 9500 406384 9512
rect 405056 9472 406384 9500
rect 405056 9460 405062 9472
rect 406378 9460 406384 9472
rect 406436 9460 406442 9512
rect 408678 9460 408684 9512
rect 408736 9500 408742 9512
rect 411162 9500 411168 9512
rect 408736 9472 411168 9500
rect 408736 9460 408742 9472
rect 411162 9460 411168 9472
rect 411220 9460 411226 9512
rect 413922 9460 413928 9512
rect 413980 9500 413986 9512
rect 419350 9500 419356 9512
rect 413980 9472 419356 9500
rect 413980 9460 413986 9472
rect 419350 9460 419356 9472
rect 419408 9460 419414 9512
rect 432046 9460 432052 9512
rect 432104 9500 432110 9512
rect 432690 9500 432696 9512
rect 432104 9472 432696 9500
rect 432104 9460 432110 9472
rect 432690 9460 432696 9472
rect 432748 9460 432754 9512
rect 447134 9460 447140 9512
rect 447192 9500 447198 9512
rect 447870 9500 447876 9512
rect 447192 9472 447876 9500
rect 447192 9460 447198 9472
rect 447870 9460 447876 9472
rect 447928 9460 447934 9512
rect 454402 9460 454408 9512
rect 454460 9500 454466 9512
rect 467190 9500 467196 9512
rect 454460 9472 467196 9500
rect 454460 9460 454466 9472
rect 467190 9460 467196 9472
rect 467248 9460 467254 9512
rect 475838 9460 475844 9512
rect 475896 9500 475902 9512
rect 504910 9500 504916 9512
rect 475896 9472 504916 9500
rect 475896 9460 475902 9472
rect 504910 9460 504916 9472
rect 504968 9460 504974 9512
rect 520182 9460 520188 9512
rect 520240 9500 520246 9512
rect 533430 9500 533436 9512
rect 520240 9472 533436 9500
rect 520240 9460 520246 9472
rect 533430 9460 533436 9472
rect 533488 9460 533494 9512
rect 316006 9404 316448 9432
rect 317966 9392 317972 9444
rect 318024 9432 318030 9444
rect 332502 9432 332508 9444
rect 318024 9404 332508 9432
rect 318024 9392 318030 9404
rect 332502 9392 332508 9404
rect 332560 9392 332566 9444
rect 333790 9392 333796 9444
rect 333848 9432 333854 9444
rect 349062 9432 349068 9444
rect 333848 9404 349068 9432
rect 333848 9392 333854 9404
rect 349062 9392 349068 9404
rect 349120 9392 349126 9444
rect 350350 9392 350356 9444
rect 350408 9432 350414 9444
rect 368290 9432 368296 9444
rect 350408 9404 368296 9432
rect 350408 9392 350414 9404
rect 368290 9392 368296 9404
rect 368348 9392 368354 9444
rect 459462 9392 459468 9444
rect 459520 9432 459526 9444
rect 476022 9432 476028 9444
rect 459520 9404 476028 9432
rect 459520 9392 459526 9404
rect 476022 9392 476028 9404
rect 476080 9392 476086 9444
rect 477862 9392 477868 9444
rect 477920 9432 477926 9444
rect 485130 9432 485136 9444
rect 477920 9404 485136 9432
rect 477920 9392 477926 9404
rect 485130 9392 485136 9404
rect 485188 9392 485194 9444
rect 487982 9392 487988 9444
rect 488040 9432 488046 9444
rect 519630 9432 519636 9444
rect 488040 9404 519636 9432
rect 488040 9392 488046 9404
rect 519630 9392 519636 9404
rect 519688 9392 519694 9444
rect 31294 9324 31300 9376
rect 31352 9364 31358 9376
rect 59354 9364 59360 9376
rect 31352 9336 59360 9364
rect 31352 9324 31358 9336
rect 59354 9324 59360 9336
rect 59412 9324 59418 9376
rect 111978 9324 111984 9376
rect 112036 9364 112042 9376
rect 115934 9364 115940 9376
rect 112036 9336 115940 9364
rect 112036 9324 112042 9336
rect 115934 9324 115940 9336
rect 115992 9324 115998 9376
rect 126882 9324 126888 9376
rect 126940 9364 126946 9376
rect 134150 9364 134156 9376
rect 126940 9336 134156 9364
rect 126940 9324 126946 9336
rect 134150 9324 134156 9336
rect 134208 9324 134214 9376
rect 142246 9324 142252 9376
rect 142304 9364 142310 9376
rect 149330 9364 149336 9376
rect 142304 9336 149336 9364
rect 142304 9324 142310 9336
rect 149330 9324 149336 9336
rect 149388 9324 149394 9376
rect 150434 9324 150440 9376
rect 150492 9364 150498 9376
rect 155402 9364 155408 9376
rect 150492 9336 155408 9364
rect 150492 9324 150498 9336
rect 155402 9324 155408 9336
rect 155460 9324 155466 9376
rect 167086 9324 167092 9376
rect 167144 9364 167150 9376
rect 170582 9364 170588 9376
rect 167144 9336 170588 9364
rect 167144 9324 167150 9336
rect 170582 9324 170588 9336
rect 170640 9324 170646 9376
rect 241054 9324 241060 9376
rect 241112 9364 241118 9376
rect 242802 9364 242808 9376
rect 241112 9336 242808 9364
rect 241112 9324 241118 9336
rect 242802 9324 242808 9336
rect 242860 9324 242866 9376
rect 260282 9324 260288 9376
rect 260340 9364 260346 9376
rect 262122 9364 262128 9376
rect 260340 9336 262128 9364
rect 260340 9324 260346 9336
rect 262122 9324 262128 9336
rect 262180 9324 262186 9376
rect 271414 9324 271420 9376
rect 271472 9364 271478 9376
rect 273162 9364 273168 9376
rect 271472 9336 273168 9364
rect 271472 9324 271478 9336
rect 273162 9324 273168 9336
rect 273220 9324 273226 9376
rect 290642 9324 290648 9376
rect 290700 9364 290706 9376
rect 292482 9364 292488 9376
rect 290700 9336 292488 9364
rect 290700 9324 290706 9336
rect 292482 9324 292488 9336
rect 292540 9324 292546 9376
rect 316034 9324 316040 9376
rect 316092 9364 316098 9376
rect 323302 9364 323308 9376
rect 316092 9336 323308 9364
rect 316092 9324 316098 9336
rect 323302 9324 323308 9336
rect 323360 9324 323366 9376
rect 323394 9324 323400 9376
rect 323452 9364 323458 9376
rect 331030 9364 331036 9376
rect 323452 9336 331036 9364
rect 323452 9324 323458 9336
rect 331030 9324 331036 9336
rect 331088 9324 331094 9376
rect 332134 9324 332140 9376
rect 332192 9364 332198 9376
rect 346578 9364 346584 9376
rect 332192 9336 346584 9364
rect 332192 9324 332198 9336
rect 346578 9324 346584 9336
rect 346636 9324 346642 9376
rect 348326 9324 348332 9376
rect 348384 9364 348390 9376
rect 368198 9364 368204 9376
rect 348384 9336 368204 9364
rect 348384 9324 348390 9336
rect 368198 9324 368204 9336
rect 368256 9324 368262 9376
rect 415118 9324 415124 9376
rect 415176 9364 415182 9376
rect 430666 9364 430672 9376
rect 415176 9336 430672 9364
rect 415176 9324 415182 9336
rect 430666 9324 430672 9336
rect 430724 9324 430730 9376
rect 463602 9324 463608 9376
rect 463660 9364 463666 9376
rect 478874 9364 478880 9376
rect 463660 9336 478880 9364
rect 463660 9324 463666 9336
rect 478874 9324 478880 9336
rect 478932 9324 478938 9376
rect 496078 9324 496084 9376
rect 496136 9364 496142 9376
rect 498010 9364 498016 9376
rect 496136 9336 498016 9364
rect 496136 9324 496142 9336
rect 498010 9324 498016 9336
rect 498068 9324 498074 9376
rect 498194 9324 498200 9376
rect 498252 9364 498258 9376
rect 536098 9364 536104 9376
rect 498252 9336 536104 9364
rect 498252 9324 498258 9336
rect 536098 9324 536104 9336
rect 536156 9324 536162 9376
rect 25314 9256 25320 9308
rect 25372 9296 25378 9308
rect 54202 9296 54208 9308
rect 25372 9268 54208 9296
rect 25372 9256 25378 9268
rect 54202 9256 54208 9268
rect 54260 9256 54266 9308
rect 132586 9256 132592 9308
rect 132644 9296 132650 9308
rect 140222 9296 140228 9308
rect 132644 9268 140228 9296
rect 132644 9256 132650 9268
rect 140222 9256 140228 9268
rect 140280 9256 140286 9308
rect 158990 9256 158996 9308
rect 159048 9296 159054 9308
rect 163498 9296 163504 9308
rect 159048 9268 163504 9296
rect 159048 9256 159054 9268
rect 163498 9256 163504 9268
rect 163556 9256 163562 9308
rect 169938 9256 169944 9308
rect 169996 9296 170002 9308
rect 172606 9296 172612 9308
rect 169996 9268 172612 9296
rect 169996 9256 170002 9268
rect 172606 9256 172612 9268
rect 172664 9256 172670 9308
rect 216858 9256 216864 9308
rect 216916 9296 216922 9308
rect 218146 9296 218152 9308
rect 216916 9268 218152 9296
rect 216916 9256 216922 9268
rect 218146 9256 218152 9268
rect 218204 9256 218210 9308
rect 249150 9256 249156 9308
rect 249208 9296 249214 9308
rect 249794 9296 249800 9308
rect 249208 9268 249800 9296
rect 249208 9256 249214 9268
rect 249794 9256 249800 9268
rect 249852 9256 249858 9308
rect 272426 9256 272432 9308
rect 272484 9296 272490 9308
rect 274450 9296 274456 9308
rect 272484 9268 274456 9296
rect 272484 9256 272490 9268
rect 274450 9256 274456 9268
rect 274508 9256 274514 9308
rect 284202 9256 284208 9308
rect 284260 9296 284266 9308
rect 285582 9296 285588 9308
rect 284260 9268 285588 9296
rect 284260 9256 284266 9268
rect 285582 9256 285588 9268
rect 285640 9256 285646 9308
rect 299382 9256 299388 9308
rect 299440 9296 299446 9308
rect 299934 9296 299940 9308
rect 299440 9268 299940 9296
rect 299440 9256 299446 9268
rect 299934 9256 299940 9268
rect 299992 9256 299998 9308
rect 308858 9256 308864 9308
rect 308916 9296 308922 9308
rect 308916 9268 319116 9296
rect 308916 9256 308922 9268
rect 19426 9188 19432 9240
rect 19484 9228 19490 9240
rect 49142 9228 49148 9240
rect 19484 9200 49148 9228
rect 19484 9188 19490 9200
rect 49142 9188 49148 9200
rect 49200 9188 49206 9240
rect 88518 9188 88524 9240
rect 88576 9228 88582 9240
rect 102778 9228 102784 9240
rect 88576 9200 102784 9228
rect 88576 9188 88582 9200
rect 102778 9188 102784 9200
rect 102836 9188 102842 9240
rect 111058 9188 111064 9240
rect 111116 9228 111122 9240
rect 117038 9228 117044 9240
rect 111116 9200 117044 9228
rect 111116 9188 111122 9200
rect 117038 9188 117044 9200
rect 117096 9188 117102 9240
rect 130378 9188 130384 9240
rect 130436 9228 130442 9240
rect 138198 9228 138204 9240
rect 130436 9200 138204 9228
rect 130436 9188 130442 9200
rect 138198 9188 138204 9200
rect 138256 9188 138262 9240
rect 140038 9188 140044 9240
rect 140096 9228 140102 9240
rect 146294 9228 146300 9240
rect 140096 9200 146300 9228
rect 140096 9188 140102 9200
rect 146294 9188 146300 9200
rect 146352 9188 146358 9240
rect 148962 9188 148968 9240
rect 149020 9228 149026 9240
rect 153378 9228 153384 9240
rect 149020 9200 153384 9228
rect 149020 9188 149026 9200
rect 153378 9188 153384 9200
rect 153436 9188 153442 9240
rect 157702 9188 157708 9240
rect 157760 9228 157766 9240
rect 161658 9228 161664 9240
rect 157760 9200 161664 9228
rect 157760 9188 157766 9200
rect 161658 9188 161664 9200
rect 161716 9188 161722 9240
rect 257982 9188 257988 9240
rect 258040 9228 258046 9240
rect 258166 9228 258172 9240
rect 258040 9200 258172 9228
rect 258040 9188 258046 9200
rect 258166 9188 258172 9200
rect 258224 9188 258230 9240
rect 298738 9188 298744 9240
rect 298796 9228 298802 9240
rect 300762 9228 300768 9240
rect 298796 9200 300768 9228
rect 298796 9188 298802 9200
rect 300762 9188 300768 9200
rect 300820 9188 300826 9240
rect 311802 9188 311808 9240
rect 311860 9228 311866 9240
rect 319088 9228 319116 9268
rect 322014 9256 322020 9308
rect 322072 9296 322078 9308
rect 335446 9296 335452 9308
rect 322072 9268 335452 9296
rect 322072 9256 322078 9268
rect 335446 9256 335452 9268
rect 335504 9256 335510 9308
rect 343634 9256 343640 9308
rect 343692 9296 343698 9308
rect 344646 9296 344652 9308
rect 343692 9268 344652 9296
rect 343692 9256 343698 9268
rect 344646 9256 344652 9268
rect 344704 9256 344710 9308
rect 347314 9256 347320 9308
rect 347372 9296 347378 9308
rect 367002 9296 367008 9308
rect 347372 9268 367008 9296
rect 347372 9256 347378 9268
rect 367002 9256 367008 9268
rect 367060 9256 367066 9308
rect 389818 9256 389824 9308
rect 389876 9296 389882 9308
rect 403066 9296 403072 9308
rect 389876 9268 403072 9296
rect 389876 9256 389882 9268
rect 403066 9256 403072 9268
rect 403124 9256 403130 9308
rect 424226 9256 424232 9308
rect 424284 9296 424290 9308
rect 445662 9296 445668 9308
rect 424284 9268 445668 9296
rect 424284 9256 424290 9268
rect 445662 9256 445668 9268
rect 445720 9256 445726 9308
rect 465718 9256 465724 9308
rect 465776 9296 465782 9308
rect 484302 9296 484308 9308
rect 465776 9268 484308 9296
rect 465776 9256 465782 9268
rect 484302 9256 484308 9268
rect 484360 9256 484366 9308
rect 485590 9256 485596 9308
rect 485648 9296 485654 9308
rect 529014 9296 529020 9308
rect 485648 9268 529020 9296
rect 485648 9256 485654 9268
rect 529014 9256 529020 9268
rect 529072 9256 529078 9308
rect 322106 9228 322112 9240
rect 311860 9200 319024 9228
rect 319088 9200 322112 9228
rect 311860 9188 311866 9200
rect 23014 9120 23020 9172
rect 23072 9160 23078 9172
rect 52454 9160 52460 9172
rect 23072 9132 52460 9160
rect 23072 9120 23078 9132
rect 52454 9120 52460 9132
rect 52512 9120 52518 9172
rect 88886 9120 88892 9172
rect 88944 9160 88950 9172
rect 103790 9160 103796 9172
rect 88944 9132 103796 9160
rect 88944 9120 88950 9132
rect 103790 9120 103796 9132
rect 103848 9120 103854 9172
rect 103974 9120 103980 9172
rect 104032 9160 104038 9172
rect 114922 9160 114928 9172
rect 104032 9132 114928 9160
rect 104032 9120 104038 9132
rect 114922 9120 114928 9132
rect 114980 9120 114986 9172
rect 127158 9120 127164 9172
rect 127216 9160 127222 9172
rect 136174 9160 136180 9172
rect 127216 9132 136180 9160
rect 127216 9120 127222 9132
rect 136174 9120 136180 9132
rect 136232 9120 136238 9172
rect 136542 9120 136548 9172
rect 136600 9160 136606 9172
rect 143534 9160 143540 9172
rect 136600 9132 143540 9160
rect 136600 9120 136606 9132
rect 143534 9120 143540 9132
rect 143592 9120 143598 9172
rect 150710 9120 150716 9172
rect 150768 9160 150774 9172
rect 156414 9160 156420 9172
rect 150768 9132 156420 9160
rect 150768 9120 150774 9132
rect 156414 9120 156420 9132
rect 156472 9120 156478 9172
rect 246114 9120 246120 9172
rect 246172 9160 246178 9172
rect 248322 9160 248328 9172
rect 246172 9132 248328 9160
rect 246172 9120 246178 9132
rect 248322 9120 248328 9132
rect 248380 9120 248386 9172
rect 282546 9120 282552 9172
rect 282604 9160 282610 9172
rect 284202 9160 284208 9172
rect 282604 9132 284208 9160
rect 282604 9120 282610 9132
rect 284202 9120 284208 9132
rect 284260 9120 284266 9172
rect 289630 9120 289636 9172
rect 289688 9160 289694 9172
rect 290826 9160 290832 9172
rect 289688 9132 290832 9160
rect 289688 9120 289694 9132
rect 290826 9120 290832 9132
rect 290884 9120 290890 9172
rect 314562 9120 314568 9172
rect 314620 9160 314626 9172
rect 318996 9160 319024 9200
rect 322106 9188 322112 9200
rect 322164 9188 322170 9240
rect 329742 9188 329748 9240
rect 329800 9228 329806 9240
rect 345198 9228 345204 9240
rect 329800 9200 345204 9228
rect 329800 9188 329806 9200
rect 345198 9188 345204 9200
rect 345256 9188 345262 9240
rect 351362 9188 351368 9240
rect 351420 9228 351426 9240
rect 365438 9228 365444 9240
rect 351420 9200 365444 9228
rect 351420 9188 351426 9200
rect 365438 9188 365444 9200
rect 365496 9188 365502 9240
rect 365530 9188 365536 9240
rect 365588 9228 365594 9240
rect 370130 9228 370136 9240
rect 365588 9200 370136 9228
rect 365588 9188 365594 9200
rect 370130 9188 370136 9200
rect 370188 9188 370194 9240
rect 371418 9188 371424 9240
rect 371476 9228 371482 9240
rect 391382 9228 391388 9240
rect 371476 9200 391388 9228
rect 371476 9188 371482 9200
rect 391382 9188 391388 9200
rect 391440 9188 391446 9240
rect 402790 9188 402796 9240
rect 402848 9228 402854 9240
rect 431954 9228 431960 9240
rect 402848 9200 431960 9228
rect 402848 9188 402854 9200
rect 431954 9188 431960 9200
rect 432012 9188 432018 9240
rect 445478 9188 445484 9240
rect 445536 9228 445542 9240
rect 464062 9228 464068 9240
rect 445536 9200 464068 9228
rect 445536 9188 445542 9200
rect 464062 9188 464068 9200
rect 464120 9188 464126 9240
rect 474642 9188 474648 9240
rect 474700 9228 474706 9240
rect 492582 9228 492588 9240
rect 474700 9200 492588 9228
rect 474700 9188 474706 9200
rect 492582 9188 492588 9200
rect 492640 9188 492646 9240
rect 503162 9188 503168 9240
rect 503220 9228 503226 9240
rect 546494 9228 546500 9240
rect 503220 9200 546500 9228
rect 503220 9188 503226 9200
rect 546494 9188 546500 9200
rect 546552 9188 546558 9240
rect 325602 9160 325608 9172
rect 314620 9132 316034 9160
rect 318996 9132 325608 9160
rect 314620 9120 314626 9132
rect 15930 9052 15936 9104
rect 15988 9092 15994 9104
rect 46106 9092 46112 9104
rect 15988 9064 46112 9092
rect 15988 9052 15994 9064
rect 46106 9052 46112 9064
rect 46164 9052 46170 9104
rect 64322 9052 64328 9104
rect 64380 9092 64386 9104
rect 87598 9092 87604 9104
rect 64380 9064 87604 9092
rect 64380 9052 64386 9064
rect 87598 9052 87604 9064
rect 87656 9052 87662 9104
rect 98546 9052 98552 9104
rect 98604 9092 98610 9104
rect 101766 9092 101772 9104
rect 98604 9064 101772 9092
rect 98604 9052 98610 9064
rect 101766 9052 101772 9064
rect 101824 9052 101830 9104
rect 103330 9052 103336 9104
rect 103388 9092 103394 9104
rect 120994 9092 121000 9104
rect 103388 9064 121000 9092
rect 103388 9052 103394 9064
rect 120994 9052 121000 9064
rect 121052 9052 121058 9104
rect 131114 9052 131120 9104
rect 131172 9092 131178 9104
rect 139394 9092 139400 9104
rect 131172 9064 139400 9092
rect 131172 9052 131178 9064
rect 139394 9052 139400 9064
rect 139452 9052 139458 9104
rect 155310 9052 155316 9104
rect 155368 9092 155374 9104
rect 159450 9092 159456 9104
rect 155368 9064 159456 9092
rect 155368 9052 155374 9064
rect 159450 9052 159456 9064
rect 159508 9052 159514 9104
rect 277302 9052 277308 9104
rect 277360 9092 277366 9104
rect 277670 9092 277676 9104
rect 277360 9064 277676 9092
rect 277360 9052 277366 9064
rect 277670 9052 277676 9064
rect 277728 9052 277734 9104
rect 316006 9092 316034 9132
rect 325602 9120 325608 9132
rect 325660 9120 325666 9172
rect 331122 9120 331128 9172
rect 331180 9160 331186 9172
rect 346486 9160 346492 9172
rect 331180 9132 346492 9160
rect 331180 9120 331186 9132
rect 346486 9120 346492 9132
rect 346544 9120 346550 9172
rect 356054 9120 356060 9172
rect 356112 9160 356118 9172
rect 377674 9160 377680 9172
rect 356112 9132 377680 9160
rect 356112 9120 356118 9132
rect 377674 9120 377680 9132
rect 377732 9120 377738 9172
rect 383562 9120 383568 9172
rect 383620 9160 383626 9172
rect 400030 9160 400036 9172
rect 383620 9132 400036 9160
rect 383620 9120 383626 9132
rect 400030 9120 400036 9132
rect 400088 9120 400094 9172
rect 419166 9120 419172 9172
rect 419224 9160 419230 9172
rect 450906 9160 450912 9172
rect 419224 9132 450912 9160
rect 419224 9120 419230 9132
rect 450906 9120 450912 9132
rect 450964 9120 450970 9172
rect 451182 9120 451188 9172
rect 451240 9160 451246 9172
rect 474090 9160 474096 9172
rect 451240 9132 474096 9160
rect 451240 9120 451246 9132
rect 474090 9120 474096 9132
rect 474148 9120 474154 9172
rect 481542 9120 481548 9172
rect 481600 9160 481606 9172
rect 498286 9160 498292 9172
rect 481600 9132 498292 9160
rect 481600 9120 481606 9132
rect 498286 9120 498292 9132
rect 498344 9120 498350 9172
rect 504174 9120 504180 9172
rect 504232 9160 504238 9172
rect 550266 9160 550272 9172
rect 504232 9132 550272 9160
rect 504232 9120 504238 9132
rect 550266 9120 550272 9132
rect 550324 9120 550330 9172
rect 327074 9092 327080 9104
rect 316006 9064 327080 9092
rect 327074 9052 327080 9064
rect 327132 9052 327138 9104
rect 327994 9052 328000 9104
rect 328052 9092 328058 9104
rect 332686 9092 332692 9104
rect 328052 9064 332692 9092
rect 328052 9052 328058 9064
rect 332686 9052 332692 9064
rect 332744 9052 332750 9104
rect 336182 9052 336188 9104
rect 336240 9092 336246 9104
rect 354030 9092 354036 9104
rect 336240 9064 354036 9092
rect 336240 9052 336246 9064
rect 354030 9052 354036 9064
rect 354088 9052 354094 9104
rect 354398 9052 354404 9104
rect 354456 9092 354462 9104
rect 375282 9092 375288 9104
rect 354456 9064 375288 9092
rect 354456 9052 354462 9064
rect 375282 9052 375288 9064
rect 375340 9052 375346 9104
rect 381722 9052 381728 9104
rect 381780 9092 381786 9104
rect 401594 9092 401600 9104
rect 381780 9064 401600 9092
rect 381780 9052 381786 9064
rect 401594 9052 401600 9064
rect 401652 9052 401658 9104
rect 405642 9052 405648 9104
rect 405700 9092 405706 9104
rect 421466 9092 421472 9104
rect 405700 9064 421472 9092
rect 405700 9052 405706 9064
rect 421466 9052 421472 9064
rect 421524 9052 421530 9104
rect 424870 9052 424876 9104
rect 424928 9092 424934 9104
rect 458082 9092 458088 9104
rect 424928 9064 458088 9092
rect 424928 9052 424934 9064
rect 458082 9052 458088 9064
rect 458140 9052 458146 9104
rect 466362 9052 466368 9104
rect 466420 9092 466426 9104
rect 495434 9092 495440 9104
rect 466420 9064 495440 9092
rect 466420 9052 466426 9064
rect 495434 9052 495440 9064
rect 495492 9052 495498 9104
rect 498102 9052 498108 9104
rect 498160 9092 498166 9104
rect 543182 9092 543188 9104
rect 498160 9064 543188 9092
rect 498160 9052 498166 9064
rect 543182 9052 543188 9064
rect 543240 9052 543246 9104
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 41046 9024 41052 9036
rect 10008 8996 41052 9024
rect 10008 8984 10014 8996
rect 41046 8984 41052 8996
rect 41104 8984 41110 9036
rect 57238 8984 57244 9036
rect 57296 9024 57302 9036
rect 81526 9024 81532 9036
rect 57296 8996 81532 9024
rect 57296 8984 57302 8996
rect 81526 8984 81532 8996
rect 81584 8984 81590 9036
rect 99834 8984 99840 9036
rect 99892 9024 99898 9036
rect 117958 9024 117964 9036
rect 99892 8996 117964 9024
rect 99892 8984 99898 8996
rect 117958 8984 117964 8996
rect 118016 8984 118022 9036
rect 133874 8984 133880 9036
rect 133932 9024 133938 9036
rect 142338 9024 142344 9036
rect 133932 8996 142344 9024
rect 133932 8984 133938 8996
rect 142338 8984 142344 8996
rect 142396 8984 142402 9036
rect 160094 8984 160100 9036
rect 160152 9024 160158 9036
rect 164510 9024 164516 9036
rect 160152 8996 164516 9024
rect 160152 8984 160158 8996
rect 164510 8984 164516 8996
rect 164568 8984 164574 9036
rect 177942 8984 177948 9036
rect 178000 9024 178006 9036
rect 178678 9024 178684 9036
rect 178000 8996 178684 9024
rect 178000 8984 178006 8996
rect 178678 8984 178684 8996
rect 178736 8984 178742 9036
rect 209774 8984 209780 9036
rect 209832 9024 209838 9036
rect 212074 9024 212080 9036
rect 209832 8996 212080 9024
rect 209832 8984 209838 8996
rect 212074 8984 212080 8996
rect 212132 8984 212138 9036
rect 268378 8984 268384 9036
rect 268436 9024 268442 9036
rect 269114 9024 269120 9036
rect 268436 8996 269120 9024
rect 268436 8984 268442 8996
rect 269114 8984 269120 8996
rect 269172 8984 269178 9036
rect 291654 8984 291660 9036
rect 291712 9024 291718 9036
rect 293770 9024 293776 9036
rect 291712 8996 293776 9024
rect 291712 8984 291718 8996
rect 293770 8984 293776 8996
rect 293828 8984 293834 9036
rect 302786 8984 302792 9036
rect 302844 9024 302850 9036
rect 304902 9024 304908 9036
rect 302844 8996 304908 9024
rect 302844 8984 302850 8996
rect 304902 8984 304908 8996
rect 304960 8984 304966 9036
rect 315850 8984 315856 9036
rect 315908 9024 315914 9036
rect 329650 9024 329656 9036
rect 315908 8996 329656 9024
rect 315908 8984 315914 8996
rect 329650 8984 329656 8996
rect 329708 8984 329714 9036
rect 346302 8984 346308 9036
rect 346360 9024 346366 9036
rect 365806 9024 365812 9036
rect 346360 8996 365812 9024
rect 346360 8984 346366 8996
rect 365806 8984 365812 8996
rect 365864 8984 365870 9036
rect 369578 8984 369584 9036
rect 369636 9024 369642 9036
rect 389726 9024 389732 9036
rect 369636 8996 389732 9024
rect 369636 8984 369642 8996
rect 389726 8984 389732 8996
rect 389784 8984 389790 9036
rect 401962 8984 401968 9036
rect 402020 9024 402026 9036
rect 418798 9024 418804 9036
rect 402020 8996 418804 9024
rect 402020 8984 402026 8996
rect 418798 8984 418804 8996
rect 418856 8984 418862 9036
rect 420822 8984 420828 9036
rect 420880 9024 420886 9036
rect 453298 9024 453304 9036
rect 420880 8996 453304 9024
rect 420880 8984 420886 8996
rect 453298 8984 453304 8996
rect 453356 8984 453362 9036
rect 467742 8984 467748 9036
rect 467800 9024 467806 9036
rect 507670 9024 507676 9036
rect 467800 8996 507676 9024
rect 467800 8984 467806 8996
rect 507670 8984 507676 8996
rect 507728 8984 507734 9036
rect 515122 8984 515128 9036
rect 515180 9024 515186 9036
rect 563238 9024 563244 9036
rect 515180 8996 563244 9024
rect 515180 8984 515186 8996
rect 563238 8984 563244 8996
rect 563296 8984 563302 9036
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 38010 8956 38016 8968
rect 6512 8928 38016 8956
rect 6512 8916 6518 8928
rect 38010 8916 38016 8928
rect 38068 8916 38074 8968
rect 50154 8916 50160 8968
rect 50212 8956 50218 8968
rect 75454 8956 75460 8968
rect 50212 8928 75460 8956
rect 50212 8916 50218 8928
rect 75454 8916 75460 8928
rect 75512 8916 75518 8968
rect 92750 8916 92756 8968
rect 92808 8956 92814 8968
rect 111794 8956 111800 8968
rect 92808 8928 111800 8956
rect 92808 8916 92814 8928
rect 111794 8916 111800 8928
rect 111852 8916 111858 8968
rect 111886 8916 111892 8968
rect 111944 8956 111950 8968
rect 123018 8956 123024 8968
rect 111944 8928 123024 8956
rect 111944 8916 111950 8928
rect 123018 8916 123024 8928
rect 123076 8916 123082 8968
rect 129642 8916 129648 8968
rect 129700 8956 129706 8968
rect 137186 8956 137192 8968
rect 129700 8928 137192 8956
rect 129700 8916 129706 8928
rect 137186 8916 137192 8928
rect 137244 8916 137250 8968
rect 138198 8916 138204 8968
rect 138256 8956 138262 8968
rect 145282 8956 145288 8968
rect 138256 8928 145288 8956
rect 138256 8916 138262 8928
rect 145282 8916 145288 8928
rect 145340 8916 145346 8968
rect 149698 8916 149704 8968
rect 149756 8956 149762 8968
rect 154574 8956 154580 8968
rect 149756 8928 154580 8956
rect 149756 8916 149762 8928
rect 154574 8916 154580 8928
rect 154632 8916 154638 8968
rect 286594 8916 286600 8968
rect 286652 8956 286658 8968
rect 287330 8956 287336 8968
rect 286652 8928 287336 8956
rect 286652 8916 286658 8928
rect 287330 8916 287336 8928
rect 287388 8916 287394 8968
rect 303430 8916 303436 8968
rect 303488 8956 303494 8968
rect 316218 8956 316224 8968
rect 303488 8928 316224 8956
rect 303488 8916 303494 8928
rect 316218 8916 316224 8928
rect 316276 8916 316282 8968
rect 316954 8916 316960 8968
rect 317012 8956 317018 8968
rect 323394 8956 323400 8968
rect 317012 8928 323400 8956
rect 317012 8916 317018 8928
rect 323394 8916 323400 8928
rect 323452 8916 323458 8968
rect 323486 8916 323492 8968
rect 323544 8956 323550 8968
rect 331214 8956 331220 8968
rect 323544 8928 331220 8956
rect 323544 8916 323550 8928
rect 331214 8916 331220 8928
rect 331272 8916 331278 8968
rect 339218 8916 339224 8968
rect 339276 8956 339282 8968
rect 356054 8956 356060 8968
rect 339276 8928 356060 8956
rect 339276 8916 339282 8928
rect 356054 8916 356060 8928
rect 356112 8916 356118 8968
rect 361482 8916 361488 8968
rect 361540 8956 361546 8968
rect 383562 8956 383568 8968
rect 361540 8928 383568 8956
rect 361540 8916 361546 8928
rect 383562 8916 383568 8928
rect 383620 8916 383626 8968
rect 390462 8916 390468 8968
rect 390520 8956 390526 8968
rect 413830 8956 413836 8968
rect 390520 8928 413836 8956
rect 390520 8916 390526 8928
rect 413830 8916 413836 8928
rect 413888 8916 413894 8968
rect 431310 8916 431316 8968
rect 431368 8956 431374 8968
rect 465166 8956 465172 8968
rect 431368 8928 465172 8956
rect 431368 8916 431374 8928
rect 465166 8916 465172 8928
rect 465224 8916 465230 8968
rect 473814 8916 473820 8968
rect 473872 8956 473878 8968
rect 514754 8956 514760 8968
rect 473872 8928 514760 8956
rect 473872 8916 473878 8928
rect 514754 8916 514760 8928
rect 514812 8916 514818 8968
rect 526070 8916 526076 8968
rect 526128 8956 526134 8968
rect 576302 8956 576308 8968
rect 526128 8928 576308 8956
rect 526128 8916 526134 8928
rect 576302 8916 576308 8928
rect 576360 8916 576366 8968
rect 142338 8848 142344 8900
rect 142396 8888 142402 8900
rect 148318 8888 148324 8900
rect 142396 8860 148324 8888
rect 142396 8848 142402 8860
rect 148318 8848 148324 8860
rect 148376 8848 148382 8900
rect 162854 8848 162860 8900
rect 162912 8888 162918 8900
rect 166534 8888 166540 8900
rect 162912 8860 166540 8888
rect 162912 8848 162918 8860
rect 166534 8848 166540 8860
rect 166592 8848 166598 8900
rect 214466 8848 214472 8900
rect 214524 8888 214530 8900
rect 216122 8888 216128 8900
rect 214524 8860 216128 8888
rect 214524 8848 214530 8860
rect 216122 8848 216128 8860
rect 216180 8848 216186 8900
rect 242710 8848 242716 8900
rect 242768 8888 242774 8900
rect 243262 8888 243268 8900
rect 242768 8860 243268 8888
rect 242768 8848 242774 8860
rect 243262 8848 243268 8860
rect 243320 8848 243326 8900
rect 255130 8848 255136 8900
rect 255188 8888 255194 8900
rect 256602 8888 256608 8900
rect 255188 8860 256608 8888
rect 255188 8848 255194 8860
rect 256602 8848 256608 8860
rect 256660 8848 256666 8900
rect 266262 8848 266268 8900
rect 266320 8888 266326 8900
rect 266722 8888 266728 8900
rect 266320 8860 266728 8888
rect 266320 8848 266326 8860
rect 266722 8848 266728 8860
rect 266780 8848 266786 8900
rect 312906 8848 312912 8900
rect 312964 8888 312970 8900
rect 326798 8888 326804 8900
rect 312964 8860 326804 8888
rect 312964 8848 312970 8860
rect 326798 8848 326804 8860
rect 326856 8848 326862 8900
rect 338022 8848 338028 8900
rect 338080 8888 338086 8900
rect 353386 8888 353392 8900
rect 338080 8860 353392 8888
rect 338080 8848 338086 8860
rect 353386 8848 353392 8860
rect 353444 8848 353450 8900
rect 355410 8848 355416 8900
rect 355468 8888 355474 8900
rect 368382 8888 368388 8900
rect 355468 8860 368388 8888
rect 355468 8848 355474 8860
rect 368382 8848 368388 8860
rect 368440 8848 368446 8900
rect 398742 8848 398748 8900
rect 398800 8888 398806 8900
rect 400858 8888 400864 8900
rect 398800 8860 400864 8888
rect 398800 8848 398806 8860
rect 400858 8848 400864 8860
rect 400916 8848 400922 8900
rect 106274 8780 106280 8832
rect 106332 8820 106338 8832
rect 109034 8820 109040 8832
rect 106332 8792 109040 8820
rect 106332 8780 106338 8792
rect 109034 8780 109040 8792
rect 109092 8780 109098 8832
rect 310882 8780 310888 8832
rect 310940 8820 310946 8832
rect 324406 8820 324412 8832
rect 310940 8792 324412 8820
rect 310940 8780 310946 8792
rect 324406 8780 324412 8792
rect 324464 8780 324470 8832
rect 325050 8780 325056 8832
rect 325108 8820 325114 8832
rect 333238 8820 333244 8832
rect 325108 8792 333244 8820
rect 325108 8780 325114 8792
rect 333238 8780 333244 8792
rect 333296 8780 333302 8832
rect 335170 8780 335176 8832
rect 335228 8820 335234 8832
rect 350534 8820 350540 8832
rect 335228 8792 350540 8820
rect 335228 8780 335234 8792
rect 350534 8780 350540 8792
rect 350592 8780 350598 8832
rect 365438 8780 365444 8832
rect 365496 8820 365502 8832
rect 371142 8820 371148 8832
rect 365496 8792 371148 8820
rect 365496 8780 365502 8792
rect 371142 8780 371148 8792
rect 371200 8780 371206 8832
rect 161566 8712 161572 8764
rect 161624 8752 161630 8764
rect 165614 8752 165620 8764
rect 161624 8724 165620 8752
rect 161624 8712 161630 8724
rect 165614 8712 165620 8724
rect 165672 8712 165678 8764
rect 172514 8712 172520 8764
rect 172572 8752 172578 8764
rect 174630 8752 174636 8764
rect 172572 8724 174636 8752
rect 172572 8712 172578 8724
rect 174630 8712 174636 8724
rect 174688 8712 174694 8764
rect 205082 8712 205088 8764
rect 205140 8752 205146 8764
rect 208026 8752 208032 8764
rect 205140 8724 208032 8752
rect 205140 8712 205146 8724
rect 208026 8712 208032 8724
rect 208084 8712 208090 8764
rect 220446 8712 220452 8764
rect 220504 8752 220510 8764
rect 221182 8752 221188 8764
rect 220504 8724 221188 8752
rect 220504 8712 220510 8724
rect 221182 8712 221188 8724
rect 221240 8712 221246 8764
rect 244090 8712 244096 8764
rect 244148 8752 244154 8764
rect 244642 8752 244648 8764
rect 244148 8724 244648 8752
rect 244148 8712 244154 8724
rect 244642 8712 244648 8724
rect 244700 8712 244706 8764
rect 253198 8712 253204 8764
rect 253256 8752 253262 8764
rect 254762 8752 254768 8764
rect 253256 8724 254768 8752
rect 253256 8712 253262 8724
rect 254762 8712 254768 8724
rect 254820 8712 254826 8764
rect 264330 8712 264336 8764
rect 264388 8752 264394 8764
rect 266262 8752 266268 8764
rect 264388 8724 266268 8752
rect 264388 8712 264394 8724
rect 266262 8712 266268 8724
rect 266320 8712 266326 8764
rect 270402 8712 270408 8764
rect 270460 8752 270466 8764
rect 271782 8752 271788 8764
rect 270460 8724 271788 8752
rect 270460 8712 270466 8724
rect 271782 8712 271788 8724
rect 271840 8712 271846 8764
rect 313918 8712 313924 8764
rect 313976 8752 313982 8764
rect 327994 8752 328000 8764
rect 313976 8724 328000 8752
rect 313976 8712 313982 8724
rect 327994 8712 328000 8724
rect 328052 8712 328058 8764
rect 337194 8712 337200 8764
rect 337252 8752 337258 8764
rect 353294 8752 353300 8764
rect 337252 8724 353300 8752
rect 337252 8712 337258 8724
rect 353294 8712 353300 8724
rect 353352 8712 353358 8764
rect 248138 8644 248144 8696
rect 248196 8684 248202 8696
rect 248506 8684 248512 8696
rect 248196 8656 248512 8684
rect 248196 8644 248202 8656
rect 248506 8644 248512 8656
rect 248564 8644 248570 8696
rect 267366 8644 267372 8696
rect 267424 8684 267430 8696
rect 267734 8684 267740 8696
rect 267424 8656 267740 8684
rect 267424 8644 267430 8656
rect 267734 8644 267740 8656
rect 267792 8644 267798 8696
rect 281442 8644 281448 8696
rect 281500 8684 281506 8696
rect 282730 8684 282736 8696
rect 281500 8656 282736 8684
rect 281500 8644 281506 8656
rect 282730 8644 282736 8656
rect 282788 8644 282794 8696
rect 318610 8644 318616 8696
rect 318668 8684 318674 8696
rect 323486 8684 323492 8696
rect 318668 8656 323492 8684
rect 318668 8644 318674 8656
rect 323486 8644 323492 8656
rect 323544 8644 323550 8696
rect 326982 8644 326988 8696
rect 327040 8684 327046 8696
rect 340782 8684 340788 8696
rect 327040 8656 340788 8684
rect 327040 8644 327046 8656
rect 340782 8644 340788 8656
rect 340840 8644 340846 8696
rect 342162 8644 342168 8696
rect 342220 8684 342226 8696
rect 358630 8684 358636 8696
rect 342220 8656 358636 8684
rect 342220 8644 342226 8656
rect 358630 8644 358636 8656
rect 358688 8644 358694 8696
rect 126238 8576 126244 8628
rect 126296 8616 126302 8628
rect 129090 8616 129096 8628
rect 126296 8588 129096 8616
rect 126296 8576 126302 8588
rect 129090 8576 129096 8588
rect 129148 8576 129154 8628
rect 242066 8576 242072 8628
rect 242124 8616 242130 8628
rect 244090 8616 244096 8628
rect 242124 8588 244096 8616
rect 242124 8576 242130 8588
rect 244090 8576 244096 8588
rect 244148 8576 244154 8628
rect 250162 8576 250168 8628
rect 250220 8616 250226 8628
rect 252462 8616 252468 8628
rect 250220 8588 252468 8616
rect 250220 8576 250226 8588
rect 252462 8576 252468 8588
rect 252520 8576 252526 8628
rect 293678 8576 293684 8628
rect 293736 8616 293742 8628
rect 295058 8616 295064 8628
rect 293736 8588 295064 8616
rect 293736 8576 293742 8588
rect 295058 8576 295064 8588
rect 295116 8576 295122 8628
rect 324038 8576 324044 8628
rect 324096 8616 324102 8628
rect 330294 8616 330300 8628
rect 324096 8588 330300 8616
rect 324096 8576 324102 8588
rect 330294 8576 330300 8588
rect 330352 8576 330358 8628
rect 333146 8576 333152 8628
rect 333204 8616 333210 8628
rect 346394 8616 346400 8628
rect 333204 8588 346400 8616
rect 333204 8576 333210 8588
rect 346394 8576 346400 8588
rect 346452 8576 346458 8628
rect 348970 8576 348976 8628
rect 349028 8616 349034 8628
rect 362218 8616 362224 8628
rect 349028 8588 362224 8616
rect 349028 8576 349034 8588
rect 362218 8576 362224 8588
rect 362276 8576 362282 8628
rect 212166 8508 212172 8560
rect 212224 8548 212230 8560
rect 214098 8548 214104 8560
rect 212224 8520 214104 8548
rect 212224 8508 212230 8520
rect 214098 8508 214104 8520
rect 214156 8508 214162 8560
rect 257246 8508 257252 8560
rect 257304 8548 257310 8560
rect 258074 8548 258080 8560
rect 257304 8520 258080 8548
rect 257304 8508 257310 8520
rect 258074 8508 258080 8520
rect 258132 8508 258138 8560
rect 276474 8508 276480 8560
rect 276532 8548 276538 8560
rect 277394 8548 277400 8560
rect 276532 8520 277400 8548
rect 276532 8508 276538 8520
rect 277394 8508 277400 8520
rect 277452 8508 277458 8560
rect 279510 8508 279516 8560
rect 279568 8548 279574 8560
rect 281442 8548 281448 8560
rect 279568 8520 281448 8548
rect 279568 8508 279574 8520
rect 281442 8508 281448 8520
rect 281500 8508 281506 8560
rect 329098 8508 329104 8560
rect 329156 8548 329162 8560
rect 341978 8548 341984 8560
rect 329156 8520 341984 8548
rect 329156 8508 329162 8520
rect 341978 8508 341984 8520
rect 342036 8508 342042 8560
rect 469398 8508 469404 8560
rect 469456 8548 469462 8560
rect 471330 8548 471336 8560
rect 469456 8520 471336 8548
rect 469456 8508 469462 8520
rect 471330 8508 471336 8520
rect 471388 8508 471394 8560
rect 207382 8440 207388 8492
rect 207440 8480 207446 8492
rect 210050 8480 210056 8492
rect 207440 8452 210056 8480
rect 207440 8440 207446 8452
rect 210050 8440 210056 8452
rect 210108 8440 210114 8492
rect 238662 8440 238668 8492
rect 238720 8480 238726 8492
rect 240042 8480 240048 8492
rect 238720 8452 240048 8480
rect 238720 8440 238726 8452
rect 240042 8440 240048 8452
rect 240100 8440 240106 8492
rect 325878 8440 325884 8492
rect 325936 8480 325942 8492
rect 334158 8480 334164 8492
rect 325936 8452 334164 8480
rect 325936 8440 325942 8452
rect 334158 8440 334164 8452
rect 334216 8440 334222 8492
rect 109770 8372 109776 8424
rect 109828 8412 109834 8424
rect 113910 8412 113916 8424
rect 109828 8384 113916 8412
rect 109828 8372 109834 8384
rect 113910 8372 113916 8384
rect 113968 8372 113974 8424
rect 168466 8372 168472 8424
rect 168524 8412 168530 8424
rect 171594 8412 171600 8424
rect 168524 8384 171600 8412
rect 168524 8372 168530 8384
rect 171594 8372 171600 8384
rect 171652 8372 171658 8424
rect 208578 8372 208584 8424
rect 208636 8412 208642 8424
rect 211154 8412 211160 8424
rect 208636 8384 211160 8412
rect 208636 8372 208642 8384
rect 211154 8372 211160 8384
rect 211212 8372 211218 8424
rect 296530 8372 296536 8424
rect 296588 8412 296594 8424
rect 297450 8412 297456 8424
rect 296588 8384 297456 8412
rect 296588 8372 296594 8384
rect 297450 8372 297456 8384
rect 297508 8372 297514 8424
rect 305822 8372 305828 8424
rect 305880 8412 305886 8424
rect 306374 8412 306380 8424
rect 305880 8384 306380 8412
rect 305880 8372 305886 8384
rect 306374 8372 306380 8384
rect 306432 8372 306438 8424
rect 359090 8372 359096 8424
rect 359148 8412 359154 8424
rect 364334 8412 364340 8424
rect 359148 8384 364340 8412
rect 359148 8372 359154 8384
rect 364334 8372 364340 8384
rect 364392 8372 364398 8424
rect 87414 8304 87420 8356
rect 87472 8344 87478 8356
rect 94682 8344 94688 8356
rect 87472 8316 94688 8344
rect 87472 8304 87478 8316
rect 94682 8304 94688 8316
rect 94740 8304 94746 8356
rect 109678 8304 109684 8356
rect 109736 8344 109742 8356
rect 113174 8344 113180 8356
rect 109736 8316 113180 8344
rect 109736 8304 109742 8316
rect 113174 8304 113180 8316
rect 113232 8304 113238 8356
rect 137094 8304 137100 8356
rect 137152 8344 137158 8356
rect 144270 8344 144276 8356
rect 137152 8316 144276 8344
rect 137152 8304 137158 8316
rect 144270 8304 144276 8316
rect 144328 8304 144334 8356
rect 146938 8304 146944 8356
rect 146996 8344 147002 8356
rect 152366 8344 152372 8356
rect 146996 8316 152372 8344
rect 146996 8304 147002 8316
rect 152366 8304 152372 8316
rect 152424 8304 152430 8356
rect 158806 8304 158812 8356
rect 158864 8344 158870 8356
rect 162486 8344 162492 8356
rect 158864 8316 162492 8344
rect 158864 8304 158870 8316
rect 162486 8304 162492 8316
rect 162544 8304 162550 8356
rect 218054 8304 218060 8356
rect 218112 8344 218118 8356
rect 219526 8344 219532 8356
rect 218112 8316 219532 8344
rect 218112 8304 218118 8316
rect 219526 8304 219532 8316
rect 219584 8304 219590 8356
rect 238018 8304 238024 8356
rect 238076 8344 238082 8356
rect 239306 8344 239312 8356
rect 238076 8316 239312 8344
rect 238076 8304 238082 8316
rect 239306 8304 239312 8316
rect 239364 8304 239370 8356
rect 295702 8304 295708 8356
rect 295760 8344 295766 8356
rect 296714 8344 296720 8356
rect 295760 8316 296720 8344
rect 295760 8304 295766 8316
rect 296714 8304 296720 8316
rect 296772 8304 296778 8356
rect 462682 8304 462688 8356
rect 462740 8344 462746 8356
rect 462740 8316 466500 8344
rect 462740 8304 462746 8316
rect 466472 8140 466500 8316
rect 492582 8168 492588 8220
rect 492640 8208 492646 8220
rect 515950 8208 515956 8220
rect 492640 8180 515956 8208
rect 492640 8168 492646 8180
rect 515950 8168 515956 8180
rect 516008 8168 516014 8220
rect 501782 8140 501788 8152
rect 466472 8112 501788 8140
rect 501782 8100 501788 8112
rect 501840 8100 501846 8152
rect 413830 8032 413836 8084
rect 413888 8072 413894 8084
rect 417878 8072 417884 8084
rect 413888 8044 417884 8072
rect 413888 8032 413894 8044
rect 417878 8032 417884 8044
rect 417936 8032 417942 8084
rect 483934 8032 483940 8084
rect 483992 8072 483998 8084
rect 526622 8072 526628 8084
rect 483992 8044 526628 8072
rect 483992 8032 483998 8044
rect 526622 8032 526628 8044
rect 526680 8032 526686 8084
rect 491018 7964 491024 8016
rect 491076 8004 491082 8016
rect 534902 8004 534908 8016
rect 491076 7976 534908 8004
rect 491076 7964 491082 7976
rect 534902 7964 534908 7976
rect 534960 7964 534966 8016
rect 400858 7896 400864 7948
rect 400916 7936 400922 7948
rect 427262 7936 427268 7948
rect 400916 7908 427268 7936
rect 400916 7896 400922 7908
rect 427262 7896 427268 7908
rect 427320 7896 427326 7948
rect 445662 7896 445668 7948
rect 445720 7936 445726 7948
rect 456886 7936 456892 7948
rect 445720 7908 456892 7936
rect 445720 7896 445726 7908
rect 456886 7896 456892 7908
rect 456944 7896 456950 7948
rect 499114 7896 499120 7948
rect 499172 7936 499178 7948
rect 544378 7936 544384 7948
rect 499172 7908 544384 7936
rect 499172 7896 499178 7908
rect 544378 7896 544384 7908
rect 544436 7896 544442 7948
rect 411070 7828 411076 7880
rect 411128 7868 411134 7880
rect 441522 7868 441528 7880
rect 411128 7840 441528 7868
rect 411128 7828 411134 7840
rect 441522 7828 441528 7840
rect 441580 7828 441586 7880
rect 450538 7828 450544 7880
rect 450596 7868 450602 7880
rect 487614 7868 487620 7880
rect 450596 7840 487620 7868
rect 450596 7828 450602 7840
rect 487614 7828 487620 7840
rect 487672 7828 487678 7880
rect 495434 7828 495440 7880
rect 495492 7868 495498 7880
rect 506474 7868 506480 7880
rect 495492 7840 506480 7868
rect 495492 7828 495498 7840
rect 506474 7828 506480 7840
rect 506532 7828 506538 7880
rect 510890 7828 510896 7880
rect 510948 7868 510954 7880
rect 558546 7868 558552 7880
rect 510948 7840 558552 7868
rect 510948 7828 510954 7840
rect 558546 7828 558552 7840
rect 558604 7828 558610 7880
rect 47854 7760 47860 7812
rect 47912 7800 47918 7812
rect 73430 7800 73436 7812
rect 47912 7772 73436 7800
rect 47912 7760 47918 7772
rect 73430 7760 73436 7772
rect 73488 7760 73494 7812
rect 377582 7760 377588 7812
rect 377640 7800 377646 7812
rect 402514 7800 402520 7812
rect 377640 7772 402520 7800
rect 377640 7760 377646 7772
rect 402514 7760 402520 7772
rect 402572 7760 402578 7812
rect 417142 7760 417148 7812
rect 417200 7800 417206 7812
rect 448606 7800 448612 7812
rect 417200 7772 448612 7800
rect 417200 7760 417206 7772
rect 448606 7760 448612 7772
rect 448664 7760 448670 7812
rect 457622 7760 457628 7812
rect 457680 7800 457686 7812
rect 495894 7800 495900 7812
rect 457680 7772 495900 7800
rect 457680 7760 457686 7772
rect 495894 7760 495900 7772
rect 495952 7760 495958 7812
rect 506198 7760 506204 7812
rect 506256 7800 506262 7812
rect 552658 7800 552664 7812
rect 506256 7772 552664 7800
rect 506256 7760 506262 7772
rect 552658 7760 552664 7772
rect 552716 7760 552722 7812
rect 30098 7692 30104 7744
rect 30156 7732 30162 7744
rect 58250 7732 58256 7744
rect 30156 7704 58256 7732
rect 30156 7692 30162 7704
rect 58250 7692 58256 7704
rect 58308 7692 58314 7744
rect 375190 7692 375196 7744
rect 375248 7732 375254 7744
rect 400122 7732 400128 7744
rect 375248 7704 400128 7732
rect 375248 7692 375254 7704
rect 400122 7692 400128 7704
rect 400180 7692 400186 7744
rect 401594 7692 401600 7744
rect 401652 7732 401658 7744
rect 407114 7732 407120 7744
rect 401652 7704 407120 7732
rect 401652 7692 401658 7704
rect 407114 7692 407120 7704
rect 407172 7692 407178 7744
rect 413094 7732 413100 7744
rect 407224 7704 413100 7732
rect 4798 7624 4804 7676
rect 4856 7664 4862 7676
rect 34974 7664 34980 7676
rect 4856 7636 34980 7664
rect 4856 7624 4862 7636
rect 34974 7624 34980 7636
rect 35032 7624 35038 7676
rect 69106 7624 69112 7676
rect 69164 7664 69170 7676
rect 91646 7664 91652 7676
rect 69164 7636 91652 7664
rect 69164 7624 69170 7636
rect 91646 7624 91652 7636
rect 91704 7624 91710 7676
rect 386414 7624 386420 7676
rect 386472 7664 386478 7676
rect 407224 7664 407252 7704
rect 413094 7692 413100 7704
rect 413152 7692 413158 7744
rect 418062 7692 418068 7744
rect 418120 7732 418126 7744
rect 449802 7732 449808 7744
rect 418120 7704 449808 7732
rect 418120 7692 418126 7704
rect 449802 7692 449808 7704
rect 449860 7692 449866 7744
rect 456610 7692 456616 7744
rect 456668 7732 456674 7744
rect 494698 7732 494704 7744
rect 456668 7704 494704 7732
rect 456668 7692 456674 7704
rect 494698 7692 494704 7704
rect 494756 7692 494762 7744
rect 505002 7692 505008 7744
rect 505060 7732 505066 7744
rect 551462 7732 551468 7744
rect 505060 7704 551468 7732
rect 505060 7692 505066 7704
rect 551462 7692 551468 7704
rect 551520 7692 551526 7744
rect 386472 7636 407252 7664
rect 386472 7624 386478 7636
rect 426250 7624 426256 7676
rect 426308 7664 426314 7676
rect 459186 7664 459192 7676
rect 426308 7636 459192 7664
rect 426308 7624 426314 7636
rect 459186 7624 459192 7636
rect 459244 7624 459250 7676
rect 471790 7624 471796 7676
rect 471848 7664 471854 7676
rect 512454 7664 512460 7676
rect 471848 7636 512460 7664
rect 471848 7624 471854 7636
rect 512454 7624 512460 7636
rect 512512 7624 512518 7676
rect 518342 7624 518348 7676
rect 518400 7664 518406 7676
rect 566826 7664 566832 7676
rect 518400 7636 566832 7664
rect 518400 7624 518406 7636
rect 566826 7624 566832 7636
rect 566884 7624 566890 7676
rect 17034 7556 17040 7608
rect 17092 7596 17098 7608
rect 47118 7596 47124 7608
rect 17092 7568 47124 7596
rect 17092 7556 17098 7568
rect 47118 7556 47124 7568
rect 47176 7556 47182 7608
rect 58434 7556 58440 7608
rect 58492 7596 58498 7608
rect 82814 7596 82820 7608
rect 58492 7568 82820 7596
rect 58492 7556 58498 7568
rect 82814 7556 82820 7568
rect 82872 7556 82878 7608
rect 370130 7556 370136 7608
rect 370188 7596 370194 7608
rect 388254 7596 388260 7608
rect 370188 7568 388260 7596
rect 370188 7556 370194 7568
rect 388254 7556 388260 7568
rect 388312 7556 388318 7608
rect 393682 7556 393688 7608
rect 393740 7596 393746 7608
rect 421374 7596 421380 7608
rect 393740 7568 421380 7596
rect 393740 7556 393746 7568
rect 421374 7556 421380 7568
rect 421432 7556 421438 7608
rect 421466 7556 421472 7608
rect 421524 7596 421530 7608
rect 435542 7596 435548 7608
rect 421524 7568 435548 7596
rect 421524 7556 421530 7568
rect 435542 7556 435548 7568
rect 435600 7556 435606 7608
rect 469858 7596 469864 7608
rect 441586 7568 469864 7596
rect 434990 7488 434996 7540
rect 435048 7528 435054 7540
rect 441586 7528 441614 7568
rect 469858 7556 469864 7568
rect 469916 7556 469922 7608
rect 478782 7556 478788 7608
rect 478840 7596 478846 7608
rect 520734 7596 520740 7608
rect 478840 7568 520740 7596
rect 478840 7556 478846 7568
rect 520734 7556 520740 7568
rect 520792 7556 520798 7608
rect 523034 7556 523040 7608
rect 523092 7596 523098 7608
rect 572714 7596 572720 7608
rect 523092 7568 572720 7596
rect 523092 7556 523098 7568
rect 572714 7556 572720 7568
rect 572772 7556 572778 7608
rect 435048 7500 441614 7528
rect 435048 7488 435054 7500
rect 555418 6808 555424 6860
rect 555476 6848 555482 6860
rect 580166 6848 580172 6860
rect 555476 6820 580172 6848
rect 555476 6808 555482 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 476022 6672 476028 6724
rect 476080 6712 476086 6724
rect 498194 6712 498200 6724
rect 476080 6684 498200 6712
rect 476080 6672 476086 6684
rect 498194 6672 498200 6684
rect 498252 6672 498258 6724
rect 498286 6672 498292 6724
rect 498344 6712 498350 6724
rect 524230 6712 524236 6724
rect 498344 6684 524236 6712
rect 498344 6672 498350 6684
rect 524230 6672 524236 6684
rect 524288 6672 524294 6724
rect 485130 6604 485136 6656
rect 485188 6644 485194 6656
rect 519538 6644 519544 6656
rect 485188 6616 519544 6644
rect 485188 6604 485194 6616
rect 519538 6604 519544 6616
rect 519596 6604 519602 6656
rect 519630 6604 519636 6656
rect 519688 6644 519694 6656
rect 531314 6644 531320 6656
rect 519688 6616 531320 6644
rect 519688 6604 519694 6616
rect 531314 6604 531320 6616
rect 531372 6604 531378 6656
rect 430666 6536 430672 6588
rect 430724 6576 430730 6588
rect 446214 6576 446220 6588
rect 430724 6548 446220 6576
rect 430724 6536 430730 6548
rect 446214 6536 446220 6548
rect 446272 6536 446278 6588
rect 498010 6536 498016 6588
rect 498068 6576 498074 6588
rect 540790 6576 540796 6588
rect 498068 6548 540796 6576
rect 498068 6536 498074 6548
rect 540790 6536 540796 6548
rect 540848 6536 540854 6588
rect 3142 6468 3148 6520
rect 3200 6508 3206 6520
rect 6178 6508 6184 6520
rect 3200 6480 6184 6508
rect 3200 6468 3206 6480
rect 6178 6468 6184 6480
rect 6236 6468 6242 6520
rect 400030 6468 400036 6520
rect 400088 6508 400094 6520
rect 409598 6508 409604 6520
rect 400088 6480 409604 6508
rect 400088 6468 400094 6480
rect 409598 6468 409604 6480
rect 409656 6468 409662 6520
rect 418798 6468 418804 6520
rect 418856 6508 418862 6520
rect 430850 6508 430856 6520
rect 418856 6480 430856 6508
rect 418856 6468 418862 6480
rect 430850 6468 430856 6480
rect 430908 6468 430914 6520
rect 440326 6468 440332 6520
rect 440384 6508 440390 6520
rect 476942 6508 476948 6520
rect 440384 6480 476948 6508
rect 440384 6468 440390 6480
rect 476942 6468 476948 6480
rect 477000 6468 477006 6520
rect 492766 6468 492772 6520
rect 492824 6508 492830 6520
rect 538398 6508 538404 6520
rect 492824 6480 538404 6508
rect 492824 6468 492830 6480
rect 538398 6468 538404 6480
rect 538456 6468 538462 6520
rect 374178 6400 374184 6452
rect 374236 6440 374242 6452
rect 398926 6440 398932 6452
rect 374236 6412 398932 6440
rect 374236 6400 374242 6412
rect 398926 6400 398932 6412
rect 398984 6400 398990 6452
rect 407206 6400 407212 6452
rect 407264 6440 407270 6452
rect 437934 6440 437940 6452
rect 407264 6412 437940 6440
rect 407264 6400 407270 6412
rect 437934 6400 437940 6412
rect 437992 6400 437998 6452
rect 447226 6400 447232 6452
rect 447284 6440 447290 6452
rect 484026 6440 484032 6452
rect 447284 6412 484032 6440
rect 447284 6400 447290 6412
rect 484026 6400 484032 6412
rect 484084 6400 484090 6452
rect 484302 6400 484308 6452
rect 484360 6440 484366 6452
rect 505370 6440 505376 6452
rect 484360 6412 505376 6440
rect 484360 6400 484366 6412
rect 505370 6400 505376 6412
rect 505428 6400 505434 6452
rect 507946 6400 507952 6452
rect 508004 6440 508010 6452
rect 554958 6440 554964 6452
rect 508004 6412 554964 6440
rect 508004 6400 508010 6412
rect 554958 6400 554964 6412
rect 555016 6400 555022 6452
rect 378226 6332 378232 6384
rect 378284 6372 378290 6384
rect 403618 6372 403624 6384
rect 378284 6344 403624 6372
rect 378284 6332 378290 6344
rect 403618 6332 403624 6344
rect 403676 6332 403682 6384
rect 411254 6332 411260 6384
rect 411312 6372 411318 6384
rect 442626 6372 442632 6384
rect 411312 6344 442632 6372
rect 411312 6332 411318 6344
rect 442626 6332 442632 6344
rect 442684 6332 442690 6384
rect 452746 6332 452752 6384
rect 452804 6372 452810 6384
rect 491110 6372 491116 6384
rect 452804 6344 491116 6372
rect 452804 6332 452810 6344
rect 491110 6332 491116 6344
rect 491168 6332 491174 6384
rect 501046 6332 501052 6384
rect 501104 6372 501110 6384
rect 547874 6372 547880 6384
rect 501104 6344 547880 6372
rect 501104 6332 501110 6344
rect 547874 6332 547880 6344
rect 547932 6332 547938 6384
rect 26510 6264 26516 6316
rect 26568 6304 26574 6316
rect 55306 6304 55312 6316
rect 26568 6276 55312 6304
rect 26568 6264 26574 6276
rect 55306 6264 55312 6276
rect 55364 6264 55370 6316
rect 76190 6264 76196 6316
rect 76248 6304 76254 6316
rect 98086 6304 98092 6316
rect 76248 6276 98092 6304
rect 76248 6264 76254 6276
rect 98086 6264 98092 6276
rect 98144 6264 98150 6316
rect 371878 6264 371884 6316
rect 371936 6304 371942 6316
rect 389450 6304 389456 6316
rect 371936 6276 389456 6304
rect 371936 6264 371942 6276
rect 389450 6264 389456 6276
rect 389508 6264 389514 6316
rect 392026 6264 392032 6316
rect 392084 6304 392090 6316
rect 419534 6304 419540 6316
rect 392084 6276 419540 6304
rect 392084 6264 392090 6276
rect 419534 6264 419540 6276
rect 419592 6264 419598 6316
rect 419626 6264 419632 6316
rect 419684 6304 419690 6316
rect 452102 6304 452108 6316
rect 419684 6276 452108 6304
rect 419684 6264 419690 6276
rect 452102 6264 452108 6276
rect 452160 6264 452166 6316
rect 459646 6264 459652 6316
rect 459704 6304 459710 6316
rect 499390 6304 499396 6316
rect 459704 6276 499396 6304
rect 459704 6264 459710 6276
rect 499390 6264 499396 6276
rect 499448 6264 499454 6316
rect 508038 6264 508044 6316
rect 508096 6304 508102 6316
rect 556154 6304 556160 6316
rect 508096 6276 556160 6304
rect 508096 6264 508102 6276
rect 556154 6264 556160 6276
rect 556212 6264 556218 6316
rect 2774 6196 2780 6248
rect 2832 6236 2838 6248
rect 33226 6236 33232 6248
rect 2832 6208 33232 6236
rect 2832 6196 2838 6208
rect 33226 6196 33232 6208
rect 33284 6196 33290 6248
rect 37182 6196 37188 6248
rect 37240 6236 37246 6248
rect 63402 6236 63408 6248
rect 37240 6208 63408 6236
rect 37240 6196 37246 6208
rect 63402 6196 63408 6208
rect 63460 6196 63466 6248
rect 65518 6196 65524 6248
rect 65576 6236 65582 6248
rect 88334 6236 88340 6248
rect 65576 6208 88340 6236
rect 65576 6196 65582 6208
rect 88334 6196 88340 6208
rect 88392 6196 88398 6248
rect 361574 6196 361580 6248
rect 361632 6236 361638 6248
rect 384758 6236 384764 6248
rect 361632 6208 384764 6236
rect 361632 6196 361638 6208
rect 384758 6196 384764 6208
rect 384816 6196 384822 6248
rect 396074 6196 396080 6248
rect 396132 6236 396138 6248
rect 396132 6208 422294 6236
rect 396132 6196 396138 6208
rect 12342 6128 12348 6180
rect 12400 6168 12406 6180
rect 42794 6168 42800 6180
rect 12400 6140 42800 6168
rect 12400 6128 12406 6140
rect 42794 6128 42800 6140
rect 42852 6128 42858 6180
rect 54938 6128 54944 6180
rect 54996 6168 55002 6180
rect 78766 6168 78772 6180
rect 54996 6140 78772 6168
rect 54996 6128 55002 6140
rect 78766 6128 78772 6140
rect 78824 6128 78830 6180
rect 352006 6128 352012 6180
rect 352064 6168 352070 6180
rect 374086 6168 374092 6180
rect 352064 6140 374092 6168
rect 352064 6128 352070 6140
rect 374086 6128 374092 6140
rect 374144 6128 374150 6180
rect 386414 6128 386420 6180
rect 386472 6168 386478 6180
rect 414290 6168 414296 6180
rect 386472 6140 414296 6168
rect 386472 6128 386478 6140
rect 414290 6128 414296 6140
rect 414348 6128 414354 6180
rect 422266 6168 422294 6208
rect 426526 6196 426532 6248
rect 426584 6236 426590 6248
rect 460382 6236 460388 6248
rect 426584 6208 460388 6236
rect 426584 6196 426590 6208
rect 460382 6196 460388 6208
rect 460440 6196 460446 6248
rect 467834 6196 467840 6248
rect 467892 6236 467898 6248
rect 508866 6236 508872 6248
rect 467892 6208 508872 6236
rect 467892 6196 467898 6208
rect 508866 6196 508872 6208
rect 508924 6196 508930 6248
rect 516134 6196 516140 6248
rect 516192 6236 516198 6248
rect 565630 6236 565636 6248
rect 516192 6208 565636 6236
rect 516192 6196 516198 6208
rect 565630 6196 565636 6208
rect 565688 6196 565694 6248
rect 424962 6168 424968 6180
rect 422266 6140 424968 6168
rect 424962 6128 424968 6140
rect 425020 6128 425026 6180
rect 427906 6128 427912 6180
rect 427964 6168 427970 6180
rect 462774 6168 462780 6180
rect 427964 6140 462780 6168
rect 427964 6128 427970 6140
rect 462774 6128 462780 6140
rect 462832 6128 462838 6180
rect 471974 6128 471980 6180
rect 472032 6168 472038 6180
rect 513558 6168 513564 6180
rect 472032 6140 513564 6168
rect 472032 6128 472038 6140
rect 513558 6128 513564 6140
rect 513616 6128 513622 6180
rect 520366 6128 520372 6180
rect 520424 6168 520430 6180
rect 570322 6168 570328 6180
rect 520424 6140 570328 6168
rect 520424 6128 520430 6140
rect 570322 6128 570328 6140
rect 570380 6128 570386 6180
rect 389726 5516 389732 5568
rect 389784 5556 389790 5568
rect 393038 5556 393044 5568
rect 389784 5528 393044 5556
rect 389784 5516 389790 5528
rect 393038 5516 393044 5528
rect 393096 5516 393102 5568
rect 419534 5516 419540 5568
rect 419592 5556 419598 5568
rect 420178 5556 420184 5568
rect 419592 5528 420184 5556
rect 419592 5516 419598 5528
rect 420178 5516 420184 5528
rect 420236 5516 420242 5568
rect 478874 5380 478880 5432
rect 478932 5420 478938 5432
rect 502978 5420 502984 5432
rect 478932 5392 502984 5420
rect 478932 5380 478938 5392
rect 502978 5380 502984 5392
rect 503036 5380 503042 5432
rect 505002 5380 505008 5432
rect 505060 5420 505066 5432
rect 517146 5420 517152 5432
rect 505060 5392 517152 5420
rect 505060 5380 505066 5392
rect 517146 5380 517152 5392
rect 517204 5380 517210 5432
rect 484394 5312 484400 5364
rect 484452 5352 484458 5364
rect 527818 5352 527824 5364
rect 484452 5324 527824 5352
rect 484452 5312 484458 5324
rect 527818 5312 527824 5324
rect 527876 5312 527882 5364
rect 480254 5244 480260 5296
rect 480312 5284 480318 5296
rect 523034 5284 523040 5296
rect 480312 5256 523040 5284
rect 480312 5244 480318 5256
rect 523034 5244 523040 5256
rect 523092 5244 523098 5296
rect 525426 5244 525432 5296
rect 525484 5284 525490 5296
rect 541986 5284 541992 5296
rect 525484 5256 541992 5284
rect 525484 5244 525490 5256
rect 541986 5244 541992 5256
rect 542044 5244 542050 5296
rect 464062 5176 464068 5228
rect 464120 5216 464126 5228
rect 481726 5216 481732 5228
rect 464120 5188 481732 5216
rect 464120 5176 464126 5188
rect 481726 5176 481732 5188
rect 481784 5176 481790 5228
rect 488626 5176 488632 5228
rect 488684 5216 488690 5228
rect 533706 5216 533712 5228
rect 488684 5188 533712 5216
rect 488684 5176 488690 5188
rect 533706 5176 533712 5188
rect 533764 5176 533770 5228
rect 419350 5108 419356 5160
rect 419408 5148 419414 5160
rect 445018 5148 445024 5160
rect 419408 5120 445024 5148
rect 419408 5108 419414 5120
rect 445018 5108 445024 5120
rect 445076 5108 445082 5160
rect 467190 5108 467196 5160
rect 467248 5148 467254 5160
rect 492306 5148 492312 5160
rect 467248 5120 492312 5148
rect 467248 5108 467254 5120
rect 492306 5108 492312 5120
rect 492364 5108 492370 5160
rect 492674 5108 492680 5160
rect 492732 5148 492738 5160
rect 537202 5148 537208 5160
rect 492732 5120 537208 5148
rect 492732 5108 492738 5120
rect 537202 5108 537208 5120
rect 537260 5108 537266 5160
rect 403066 5040 403072 5092
rect 403124 5080 403130 5092
rect 416682 5080 416688 5092
rect 403124 5052 416688 5080
rect 403124 5040 403130 5052
rect 416682 5040 416688 5052
rect 416740 5040 416746 5092
rect 432138 5040 432144 5092
rect 432196 5080 432202 5092
rect 466270 5080 466276 5092
rect 432196 5052 466276 5080
rect 432196 5040 432202 5052
rect 466270 5040 466276 5052
rect 466328 5040 466334 5092
rect 485774 5040 485780 5092
rect 485832 5080 485838 5092
rect 530118 5080 530124 5092
rect 485832 5052 530124 5080
rect 485832 5040 485838 5052
rect 530118 5040 530124 5052
rect 530176 5040 530182 5092
rect 533430 5040 533436 5092
rect 533488 5080 533494 5092
rect 569126 5080 569132 5092
rect 533488 5052 569132 5080
rect 533488 5040 533494 5052
rect 569126 5040 569132 5052
rect 569184 5040 569190 5092
rect 72602 4972 72608 5024
rect 72660 5012 72666 5024
rect 87414 5012 87420 5024
rect 72660 4984 87420 5012
rect 72660 4972 72666 4984
rect 87414 4972 87420 4984
rect 87472 4972 87478 5024
rect 371234 4972 371240 5024
rect 371292 5012 371298 5024
rect 396534 5012 396540 5024
rect 371292 4984 396540 5012
rect 371292 4972 371298 4984
rect 396534 4972 396540 4984
rect 396592 4972 396598 5024
rect 406378 4972 406384 5024
rect 406436 5012 406442 5024
rect 434438 5012 434444 5024
rect 406436 4984 434444 5012
rect 406436 4972 406442 4984
rect 434438 4972 434444 4984
rect 434496 4972 434502 5024
rect 437474 4972 437480 5024
rect 437532 5012 437538 5024
rect 473446 5012 473452 5024
rect 437532 4984 473452 5012
rect 437532 4972 437538 4984
rect 473446 4972 473452 4984
rect 473504 4972 473510 5024
rect 474090 4972 474096 5024
rect 474148 5012 474154 5024
rect 488810 5012 488816 5024
rect 474148 4984 488816 5012
rect 474148 4972 474154 4984
rect 488810 4972 488816 4984
rect 488868 4972 488874 5024
rect 499666 4972 499672 5024
rect 499724 5012 499730 5024
rect 545482 5012 545488 5024
rect 499724 4984 545488 5012
rect 499724 4972 499730 4984
rect 545482 4972 545488 4984
rect 545540 4972 545546 5024
rect 21818 4904 21824 4956
rect 21876 4944 21882 4956
rect 51074 4944 51080 4956
rect 21876 4916 51080 4944
rect 21876 4904 21882 4916
rect 51074 4904 51080 4916
rect 51132 4904 51138 4956
rect 51350 4904 51356 4956
rect 51408 4944 51414 4956
rect 75914 4944 75920 4956
rect 51408 4916 75920 4944
rect 51408 4904 51414 4916
rect 75914 4904 75920 4916
rect 75972 4904 75978 4956
rect 364334 4904 364340 4956
rect 364392 4944 364398 4956
rect 381170 4944 381176 4956
rect 364392 4916 381176 4944
rect 364392 4904 364398 4916
rect 381170 4904 381176 4916
rect 381228 4904 381234 4956
rect 383654 4904 383660 4956
rect 383712 4944 383718 4956
rect 410794 4944 410800 4956
rect 383712 4916 410800 4944
rect 383712 4904 383718 4916
rect 410794 4904 410800 4916
rect 410852 4904 410858 4956
rect 411162 4904 411168 4956
rect 411220 4944 411226 4956
rect 439130 4944 439136 4956
rect 411220 4916 439136 4944
rect 411220 4904 411226 4916
rect 439130 4904 439136 4916
rect 439188 4904 439194 4956
rect 443086 4904 443092 4956
rect 443144 4944 443150 4956
rect 480530 4944 480536 4956
rect 443144 4916 480536 4944
rect 443144 4904 443150 4916
rect 480530 4904 480536 4916
rect 480588 4904 480594 4956
rect 513374 4904 513380 4956
rect 513432 4944 513438 4956
rect 562042 4944 562048 4956
rect 513432 4916 562048 4944
rect 513432 4904 513438 4916
rect 562042 4904 562048 4916
rect 562100 4904 562106 4956
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 33134 4876 33140 4888
rect 1728 4848 33140 4876
rect 1728 4836 1734 4848
rect 33134 4836 33140 4848
rect 33192 4836 33198 4888
rect 33594 4836 33600 4888
rect 33652 4876 33658 4888
rect 60734 4876 60740 4888
rect 33652 4848 60740 4876
rect 33652 4836 33658 4848
rect 60734 4836 60740 4848
rect 60792 4836 60798 4888
rect 62022 4836 62028 4888
rect 62080 4876 62086 4888
rect 85666 4876 85672 4888
rect 62080 4848 85672 4876
rect 62080 4836 62086 4848
rect 85666 4836 85672 4848
rect 85724 4836 85730 4888
rect 367278 4836 367284 4888
rect 367336 4876 367342 4888
rect 391842 4876 391848 4888
rect 367336 4848 391848 4876
rect 367336 4836 367342 4848
rect 391842 4836 391848 4848
rect 391900 4836 391906 4888
rect 394694 4836 394700 4888
rect 394752 4876 394758 4888
rect 423766 4876 423772 4888
rect 394752 4848 423772 4876
rect 394752 4836 394758 4848
rect 423766 4836 423772 4848
rect 423824 4836 423830 4888
rect 447134 4836 447140 4888
rect 447192 4876 447198 4888
rect 485222 4876 485228 4888
rect 447192 4848 485228 4876
rect 447192 4836 447198 4848
rect 485222 4836 485228 4848
rect 485280 4836 485286 4888
rect 510614 4836 510620 4888
rect 510672 4876 510678 4888
rect 559742 4876 559748 4888
rect 510672 4848 559748 4876
rect 510672 4836 510678 4848
rect 559742 4836 559748 4848
rect 559800 4836 559806 4888
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 38654 4808 38660 4820
rect 7708 4780 38660 4808
rect 7708 4768 7714 4780
rect 38654 4768 38660 4780
rect 38712 4768 38718 4820
rect 40678 4768 40684 4820
rect 40736 4808 40742 4820
rect 67726 4808 67732 4820
rect 40736 4780 67732 4808
rect 40736 4768 40742 4780
rect 67726 4768 67732 4780
rect 67784 4768 67790 4820
rect 79686 4768 79692 4820
rect 79744 4808 79750 4820
rect 100754 4808 100760 4820
rect 79744 4780 100760 4808
rect 79744 4768 79750 4780
rect 100754 4768 100760 4780
rect 100812 4768 100818 4820
rect 379514 4768 379520 4820
rect 379572 4808 379578 4820
rect 406010 4808 406016 4820
rect 379572 4780 406016 4808
rect 379572 4768 379578 4780
rect 406010 4768 406016 4780
rect 406068 4768 406074 4820
rect 422294 4768 422300 4820
rect 422352 4808 422358 4820
rect 455690 4808 455696 4820
rect 422352 4780 455696 4808
rect 422352 4768 422358 4780
rect 455690 4768 455696 4780
rect 455748 4768 455754 4820
rect 471330 4768 471336 4820
rect 471388 4808 471394 4820
rect 510062 4808 510068 4820
rect 471388 4780 510068 4808
rect 471388 4768 471394 4780
rect 510062 4768 510068 4780
rect 510120 4768 510126 4820
rect 523126 4768 523132 4820
rect 523184 4808 523190 4820
rect 573910 4808 573916 4820
rect 523184 4780 573916 4808
rect 523184 4768 523190 4780
rect 573910 4768 573916 4780
rect 573968 4768 573974 4820
rect 546494 4632 546500 4684
rect 546552 4672 546558 4684
rect 549070 4672 549076 4684
rect 546552 4644 549076 4672
rect 546552 4632 546558 4644
rect 549070 4632 549076 4644
rect 549128 4632 549134 4684
rect 391382 4292 391388 4344
rect 391440 4332 391446 4344
rect 395338 4332 395344 4344
rect 391440 4304 395344 4332
rect 391440 4292 391446 4304
rect 395338 4292 395344 4304
rect 395396 4292 395402 4344
rect 34790 4088 34796 4140
rect 34848 4128 34854 4140
rect 62114 4128 62120 4140
rect 34848 4100 62120 4128
rect 34848 4088 34854 4100
rect 62114 4088 62120 4100
rect 62172 4088 62178 4140
rect 63218 4088 63224 4140
rect 63276 4128 63282 4140
rect 85574 4128 85580 4140
rect 63276 4100 85580 4128
rect 63276 4088 63282 4100
rect 85574 4088 85580 4100
rect 85632 4088 85638 4140
rect 89162 4088 89168 4140
rect 89220 4128 89226 4140
rect 106274 4128 106280 4140
rect 89220 4100 106280 4128
rect 89220 4088 89226 4100
rect 106274 4088 106280 4100
rect 106332 4088 106338 4140
rect 116394 4088 116400 4140
rect 116452 4128 116458 4140
rect 131022 4128 131028 4140
rect 116452 4100 131028 4128
rect 116452 4088 116458 4100
rect 131022 4088 131028 4100
rect 131080 4088 131086 4140
rect 131758 4088 131764 4140
rect 131816 4128 131822 4140
rect 138198 4128 138204 4140
rect 131816 4100 138204 4128
rect 131816 4088 131822 4100
rect 138198 4088 138204 4100
rect 138256 4088 138262 4140
rect 164878 4088 164884 4140
rect 164936 4128 164942 4140
rect 171226 4128 171232 4140
rect 164936 4100 171232 4128
rect 164936 4088 164942 4100
rect 171226 4088 171232 4100
rect 171284 4088 171290 4140
rect 197906 4088 197912 4140
rect 197964 4128 197970 4140
rect 201586 4128 201592 4140
rect 197964 4100 201592 4128
rect 197964 4088 197970 4100
rect 201586 4088 201592 4100
rect 201644 4088 201650 4140
rect 247862 4088 247868 4140
rect 247920 4128 247926 4140
rect 249978 4128 249984 4140
rect 247920 4100 249984 4128
rect 247920 4088 247926 4100
rect 249978 4088 249984 4100
rect 250036 4088 250042 4140
rect 274450 4088 274456 4140
rect 274508 4128 274514 4140
rect 279510 4128 279516 4140
rect 274508 4100 279516 4128
rect 274508 4088 274514 4100
rect 279510 4088 279516 4100
rect 279568 4088 279574 4140
rect 281442 4088 281448 4140
rect 281500 4128 281506 4140
rect 287790 4128 287796 4140
rect 281500 4100 287796 4128
rect 281500 4088 281506 4100
rect 287790 4088 287796 4100
rect 287848 4088 287854 4140
rect 300762 4088 300768 4140
rect 300820 4128 300826 4140
rect 310238 4128 310244 4140
rect 300820 4100 310244 4128
rect 300820 4088 300826 4100
rect 310238 4088 310244 4100
rect 310296 4088 310302 4140
rect 362954 4088 362960 4140
rect 363012 4128 363018 4140
rect 385954 4128 385960 4140
rect 363012 4100 385960 4128
rect 363012 4088 363018 4100
rect 385954 4088 385960 4100
rect 386012 4088 386018 4140
rect 390554 4088 390560 4140
rect 390612 4128 390618 4140
rect 418982 4128 418988 4140
rect 390612 4100 418988 4128
rect 390612 4088 390618 4100
rect 418982 4088 418988 4100
rect 419040 4088 419046 4140
rect 442994 4088 443000 4140
rect 443052 4128 443058 4140
rect 479334 4128 479340 4140
rect 443052 4100 479340 4128
rect 443052 4088 443058 4100
rect 479334 4088 479340 4100
rect 479392 4088 479398 4140
rect 499574 4088 499580 4140
rect 499632 4128 499638 4140
rect 546678 4128 546684 4140
rect 499632 4100 546684 4128
rect 499632 4088 499638 4100
rect 546678 4088 546684 4100
rect 546736 4088 546742 4140
rect 24210 4020 24216 4072
rect 24268 4060 24274 4072
rect 52546 4060 52552 4072
rect 24268 4032 52552 4060
rect 24268 4020 24274 4032
rect 52546 4020 52552 4032
rect 52604 4020 52610 4072
rect 56042 4020 56048 4072
rect 56100 4060 56106 4072
rect 80054 4060 80060 4072
rect 56100 4032 80060 4060
rect 56100 4020 56106 4032
rect 80054 4020 80060 4032
rect 80112 4020 80118 4072
rect 85666 4020 85672 4072
rect 85724 4060 85730 4072
rect 105814 4060 105820 4072
rect 85724 4032 105820 4060
rect 85724 4020 85730 4032
rect 105814 4020 105820 4032
rect 105872 4020 105878 4072
rect 117590 4020 117596 4072
rect 117648 4060 117654 4072
rect 132494 4060 132500 4072
rect 117648 4032 132500 4060
rect 117648 4020 117654 4032
rect 132494 4020 132500 4032
rect 132552 4020 132558 4072
rect 136450 4020 136456 4072
rect 136508 4060 136514 4072
rect 142246 4060 142252 4072
rect 136508 4032 142252 4060
rect 136508 4020 136514 4032
rect 142246 4020 142252 4032
rect 142304 4020 142310 4072
rect 147122 4020 147128 4072
rect 147180 4060 147186 4072
rect 153194 4060 153200 4072
rect 147180 4032 153200 4060
rect 147180 4020 147186 4032
rect 153194 4020 153200 4032
rect 153252 4020 153258 4072
rect 282822 4020 282828 4072
rect 282880 4060 282886 4072
rect 288986 4060 288992 4072
rect 282880 4032 288992 4060
rect 282880 4020 282886 4032
rect 288986 4020 288992 4032
rect 289044 4020 289050 4072
rect 296714 4020 296720 4072
rect 296772 4060 296778 4072
rect 306742 4060 306748 4072
rect 296772 4032 306748 4060
rect 296772 4020 296778 4032
rect 306742 4020 306748 4032
rect 306800 4020 306806 4072
rect 394234 4060 394240 4072
rect 373966 4032 394240 4060
rect 28902 3952 28908 4004
rect 28960 3992 28966 4004
rect 56686 3992 56692 4004
rect 28960 3964 56692 3992
rect 28960 3952 28966 3964
rect 56686 3952 56692 3964
rect 56744 3952 56750 4004
rect 60826 3952 60832 4004
rect 60884 3992 60890 4004
rect 84194 3992 84200 4004
rect 60884 3964 84200 3992
rect 60884 3952 60890 3964
rect 84194 3952 84200 3964
rect 84252 3952 84258 4004
rect 86862 3952 86868 4004
rect 86920 3992 86926 4004
rect 106826 3992 106832 4004
rect 86920 3964 106832 3992
rect 86920 3952 86926 3964
rect 106826 3952 106832 3964
rect 106884 3952 106890 4004
rect 108114 3952 108120 4004
rect 108172 3992 108178 4004
rect 124306 3992 124312 4004
rect 108172 3964 124312 3992
rect 108172 3952 108178 3964
rect 124306 3952 124312 3964
rect 124364 3952 124370 4004
rect 128170 3952 128176 4004
rect 128228 3992 128234 4004
rect 133874 3992 133880 4004
rect 128228 3964 133880 3992
rect 128228 3952 128234 3964
rect 133874 3952 133880 3964
rect 133932 3952 133938 4004
rect 137646 3952 137652 4004
rect 137704 3992 137710 4004
rect 143626 3992 143632 4004
rect 137704 3964 143632 3992
rect 137704 3952 137710 3964
rect 143626 3952 143632 3964
rect 143684 3952 143690 4004
rect 166074 3952 166080 4004
rect 166132 3992 166138 4004
rect 172514 3992 172520 4004
rect 166132 3964 172520 3992
rect 166132 3952 166138 3964
rect 172514 3952 172520 3964
rect 172572 3952 172578 4004
rect 184934 3952 184940 4004
rect 184992 3992 184998 4004
rect 190454 3992 190460 4004
rect 184992 3964 190460 3992
rect 184992 3952 184998 3964
rect 190454 3952 190460 3964
rect 190512 3952 190518 4004
rect 195606 3952 195612 4004
rect 195664 3992 195670 4004
rect 200206 3992 200212 4004
rect 195664 3964 200212 3992
rect 195664 3952 195670 3964
rect 200206 3952 200212 3964
rect 200264 3952 200270 4004
rect 255222 3952 255228 4004
rect 255280 3992 255286 4004
rect 258258 3992 258264 4004
rect 255280 3964 258264 3992
rect 255280 3952 255286 3964
rect 258258 3952 258264 3964
rect 258316 3952 258322 4004
rect 273162 3952 273168 4004
rect 273220 3992 273226 4004
rect 278314 3992 278320 4004
rect 273220 3964 278320 3992
rect 273220 3952 273226 3964
rect 278314 3952 278320 3964
rect 278372 3952 278378 4004
rect 295886 3952 295892 4004
rect 295944 3992 295950 4004
rect 305546 3992 305552 4004
rect 295944 3964 305552 3992
rect 295944 3952 295950 3964
rect 305546 3952 305552 3964
rect 305604 3952 305610 4004
rect 362218 3952 362224 4004
rect 362276 3992 362282 4004
rect 369394 3992 369400 4004
rect 362276 3964 369400 3992
rect 362276 3952 362282 3964
rect 369394 3952 369400 3964
rect 369452 3952 369458 4004
rect 369854 3952 369860 4004
rect 369912 3992 369918 4004
rect 373966 3992 373994 4032
rect 394234 4020 394240 4032
rect 394292 4020 394298 4072
rect 402974 4020 402980 4072
rect 403032 4060 403038 4072
rect 433242 4060 433248 4072
rect 403032 4032 433248 4060
rect 403032 4020 403038 4032
rect 433242 4020 433248 4032
rect 433300 4020 433306 4072
rect 445754 4020 445760 4072
rect 445812 4060 445818 4072
rect 482830 4060 482836 4072
rect 445812 4032 482836 4060
rect 445812 4020 445818 4032
rect 482830 4020 482836 4032
rect 482888 4020 482894 4072
rect 518894 4020 518900 4072
rect 518952 4060 518958 4072
rect 568022 4060 568028 4072
rect 518952 4032 568028 4060
rect 518952 4020 518958 4032
rect 568022 4020 568028 4032
rect 568080 4020 568086 4072
rect 369912 3964 373994 3992
rect 369912 3952 369918 3964
rect 375374 3952 375380 4004
rect 375432 3992 375438 4004
rect 375432 3964 379008 3992
rect 375432 3952 375438 3964
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 41414 3924 41420 3936
rect 11204 3896 41420 3924
rect 11204 3884 11210 3896
rect 41414 3884 41420 3896
rect 41472 3884 41478 3936
rect 41874 3884 41880 3936
rect 41932 3924 41938 3936
rect 67634 3924 67640 3936
rect 41932 3896 67640 3924
rect 41932 3884 41938 3896
rect 67634 3884 67640 3896
rect 67692 3884 67698 3936
rect 67910 3884 67916 3936
rect 67968 3924 67974 3936
rect 89714 3924 89720 3936
rect 67968 3896 89720 3924
rect 67968 3884 67974 3896
rect 89714 3884 89720 3896
rect 89772 3884 89778 3936
rect 90358 3884 90364 3936
rect 90416 3924 90422 3936
rect 107654 3924 107660 3936
rect 90416 3896 107660 3924
rect 90416 3884 90422 3896
rect 107654 3884 107660 3896
rect 107712 3884 107718 3936
rect 110506 3884 110512 3936
rect 110564 3924 110570 3936
rect 126974 3924 126980 3936
rect 110564 3896 126980 3924
rect 110564 3884 110570 3896
rect 126974 3884 126980 3896
rect 127032 3884 127038 3936
rect 135254 3884 135260 3936
rect 135312 3924 135318 3936
rect 142338 3924 142344 3936
rect 135312 3896 142344 3924
rect 135312 3884 135318 3896
rect 142338 3884 142344 3896
rect 142396 3884 142402 3936
rect 179046 3884 179052 3936
rect 179104 3924 179110 3936
rect 185118 3924 185124 3936
rect 179104 3896 185124 3924
rect 179104 3884 179110 3896
rect 185118 3884 185124 3896
rect 185176 3884 185182 3936
rect 285582 3884 285588 3936
rect 285640 3924 285646 3936
rect 293678 3924 293684 3936
rect 285640 3896 293684 3924
rect 285640 3884 285646 3896
rect 293678 3884 293684 3896
rect 293736 3884 293742 3936
rect 299934 3884 299940 3936
rect 299992 3924 299998 3936
rect 311434 3924 311440 3936
rect 299992 3896 311440 3924
rect 299992 3884 299998 3896
rect 311434 3884 311440 3896
rect 311492 3884 311498 3936
rect 356146 3884 356152 3936
rect 356204 3924 356210 3936
rect 378870 3924 378876 3936
rect 356204 3896 378876 3924
rect 356204 3884 356210 3896
rect 378870 3884 378876 3896
rect 378928 3884 378934 3936
rect 378980 3924 379008 3964
rect 382366 3952 382372 4004
rect 382424 3992 382430 4004
rect 408402 3992 408408 4004
rect 382424 3964 408408 3992
rect 382424 3952 382430 3964
rect 408402 3952 408408 3964
rect 408460 3952 408466 4004
rect 412726 3952 412732 4004
rect 412784 3992 412790 4004
rect 443822 3992 443828 4004
rect 412784 3964 443828 3992
rect 412784 3952 412790 3964
rect 443822 3952 443828 3964
rect 443880 3952 443886 4004
rect 448514 3952 448520 4004
rect 448572 3992 448578 4004
rect 486418 3992 486424 4004
rect 448572 3964 486424 3992
rect 448572 3952 448578 3964
rect 486418 3952 486424 3964
rect 486476 3952 486482 4004
rect 511994 3952 512000 4004
rect 512052 3992 512058 4004
rect 560846 3992 560852 4004
rect 512052 3964 560852 3992
rect 512052 3952 512058 3964
rect 560846 3952 560852 3964
rect 560904 3952 560910 4004
rect 378980 3896 383654 3924
rect 18230 3816 18236 3868
rect 18288 3856 18294 3868
rect 48498 3856 48504 3868
rect 18288 3828 48504 3856
rect 18288 3816 18294 3828
rect 48498 3816 48504 3828
rect 48556 3816 48562 3868
rect 87966 3816 87972 3868
rect 88024 3856 88030 3868
rect 101950 3856 101956 3868
rect 88024 3828 101956 3856
rect 88024 3816 88030 3828
rect 101950 3816 101956 3828
rect 102008 3816 102014 3868
rect 102042 3816 102048 3868
rect 102100 3856 102106 3868
rect 104894 3856 104900 3868
rect 102100 3828 104900 3856
rect 102100 3816 102106 3828
rect 104894 3816 104900 3828
rect 104952 3816 104958 3868
rect 109310 3816 109316 3868
rect 109368 3856 109374 3868
rect 125594 3856 125600 3868
rect 109368 3828 125600 3856
rect 109368 3816 109374 3828
rect 125594 3816 125600 3828
rect 125652 3816 125658 3868
rect 125870 3816 125876 3868
rect 125928 3856 125934 3868
rect 132586 3856 132592 3868
rect 125928 3828 132592 3856
rect 125928 3816 125934 3828
rect 132586 3816 132592 3828
rect 132644 3816 132650 3868
rect 132954 3816 132960 3868
rect 133012 3856 133018 3868
rect 140038 3856 140044 3868
rect 133012 3828 140044 3856
rect 133012 3816 133018 3828
rect 140038 3816 140044 3828
rect 140096 3816 140102 3868
rect 141234 3816 141240 3868
rect 141292 3856 141298 3868
rect 148962 3856 148968 3868
rect 141292 3828 148968 3856
rect 141292 3816 141298 3828
rect 148962 3816 148968 3828
rect 149020 3816 149026 3868
rect 150618 3816 150624 3868
rect 150676 3856 150682 3868
rect 157702 3856 157708 3868
rect 150676 3828 157708 3856
rect 150676 3816 150682 3828
rect 157702 3816 157708 3828
rect 157760 3816 157766 3868
rect 161290 3816 161296 3868
rect 161348 3856 161354 3868
rect 167086 3856 167092 3868
rect 161348 3828 167092 3856
rect 161348 3816 161354 3828
rect 167086 3816 167092 3828
rect 167144 3816 167150 3868
rect 168374 3816 168380 3868
rect 168432 3856 168438 3868
rect 176562 3856 176568 3868
rect 168432 3828 176568 3856
rect 168432 3816 168438 3828
rect 176562 3816 176568 3828
rect 176620 3816 176626 3868
rect 176654 3816 176660 3868
rect 176712 3856 176718 3868
rect 183554 3856 183560 3868
rect 176712 3828 183560 3856
rect 176712 3816 176718 3828
rect 183554 3816 183560 3828
rect 183612 3816 183618 3868
rect 257890 3816 257896 3868
rect 257948 3856 257954 3868
rect 260650 3856 260656 3868
rect 257948 3828 260656 3856
rect 257948 3816 257954 3828
rect 260650 3816 260656 3828
rect 260708 3816 260714 3868
rect 264882 3816 264888 3868
rect 264940 3856 264946 3868
rect 268838 3856 268844 3868
rect 264940 3828 268844 3856
rect 264940 3816 264946 3828
rect 268838 3816 268844 3828
rect 268896 3816 268902 3868
rect 284202 3816 284208 3868
rect 284260 3856 284266 3868
rect 291378 3856 291384 3868
rect 284260 3828 291384 3856
rect 284260 3816 284266 3828
rect 291378 3816 291384 3828
rect 291436 3816 291442 3868
rect 292482 3816 292488 3868
rect 292540 3856 292546 3868
rect 300762 3856 300768 3868
rect 292540 3828 300768 3856
rect 292540 3816 292546 3828
rect 300762 3816 300768 3828
rect 300820 3816 300826 3868
rect 309042 3856 309048 3868
rect 300872 3828 309048 3856
rect 14734 3748 14740 3800
rect 14792 3788 14798 3800
rect 44174 3788 44180 3800
rect 14792 3760 44180 3788
rect 14792 3748 14798 3760
rect 44174 3748 44180 3760
rect 44232 3748 44238 3800
rect 44266 3748 44272 3800
rect 44324 3788 44330 3800
rect 70486 3788 70492 3800
rect 44324 3760 70492 3788
rect 44324 3748 44330 3760
rect 70486 3748 70492 3760
rect 70544 3748 70550 3800
rect 74994 3748 75000 3800
rect 75052 3788 75058 3800
rect 96614 3788 96620 3800
rect 75052 3760 96620 3788
rect 75052 3748 75058 3760
rect 96614 3748 96620 3760
rect 96672 3748 96678 3800
rect 97442 3748 97448 3800
rect 97500 3788 97506 3800
rect 111978 3788 111984 3800
rect 97500 3760 111984 3788
rect 97500 3748 97506 3760
rect 111978 3748 111984 3760
rect 112036 3748 112042 3800
rect 115198 3748 115204 3800
rect 115256 3788 115262 3800
rect 131298 3788 131304 3800
rect 115256 3760 131304 3788
rect 115256 3748 115262 3760
rect 131298 3748 131304 3760
rect 131356 3748 131362 3800
rect 138842 3748 138848 3800
rect 138900 3788 138906 3800
rect 146202 3788 146208 3800
rect 138900 3760 146208 3788
rect 138900 3748 138906 3760
rect 146202 3748 146208 3760
rect 146260 3748 146266 3800
rect 148318 3748 148324 3800
rect 148376 3788 148382 3800
rect 155310 3788 155316 3800
rect 148376 3760 155316 3788
rect 148376 3748 148382 3760
rect 155310 3748 155316 3760
rect 155368 3748 155374 3800
rect 158898 3748 158904 3800
rect 158956 3788 158962 3800
rect 165982 3788 165988 3800
rect 158956 3760 165988 3788
rect 158956 3748 158962 3760
rect 165982 3748 165988 3760
rect 166040 3748 166046 3800
rect 167178 3748 167184 3800
rect 167236 3788 167242 3800
rect 175182 3788 175188 3800
rect 167236 3760 175188 3788
rect 167236 3748 167242 3760
rect 175182 3748 175188 3760
rect 175240 3748 175246 3800
rect 196802 3748 196808 3800
rect 196860 3788 196866 3800
rect 200114 3788 200120 3800
rect 196860 3760 200120 3788
rect 196860 3748 196866 3760
rect 200114 3748 200120 3760
rect 200172 3748 200178 3800
rect 267642 3748 267648 3800
rect 267700 3788 267706 3800
rect 271230 3788 271236 3800
rect 267700 3760 271236 3788
rect 267700 3748 267706 3760
rect 271230 3748 271236 3760
rect 271288 3748 271294 3800
rect 274542 3748 274548 3800
rect 274600 3788 274606 3800
rect 280706 3788 280712 3800
rect 274600 3760 280712 3788
rect 274600 3748 274606 3760
rect 280706 3748 280712 3760
rect 280764 3748 280770 3800
rect 298094 3748 298100 3800
rect 298152 3788 298158 3800
rect 300872 3788 300900 3828
rect 309042 3816 309048 3828
rect 309100 3816 309106 3868
rect 341978 3816 341984 3868
rect 342036 3856 342042 3868
rect 345750 3856 345756 3868
rect 342036 3828 345756 3856
rect 342036 3816 342042 3828
rect 345750 3816 345756 3828
rect 345808 3816 345814 3868
rect 351914 3816 351920 3868
rect 351972 3856 351978 3868
rect 372890 3856 372896 3868
rect 351972 3828 372896 3856
rect 351972 3816 351978 3828
rect 372890 3816 372896 3828
rect 372948 3816 372954 3868
rect 383626 3856 383654 3896
rect 387794 3884 387800 3936
rect 387852 3924 387858 3936
rect 415486 3924 415492 3936
rect 387852 3896 415492 3924
rect 387852 3884 387858 3896
rect 415486 3884 415492 3896
rect 415544 3884 415550 3936
rect 421006 3884 421012 3936
rect 421064 3924 421070 3936
rect 454494 3924 454500 3936
rect 421064 3896 454500 3924
rect 421064 3884 421070 3896
rect 454494 3884 454500 3896
rect 454552 3884 454558 3936
rect 460934 3884 460940 3936
rect 460992 3924 460998 3936
rect 500586 3924 500592 3936
rect 460992 3896 500592 3924
rect 460992 3884 460998 3896
rect 500586 3884 500592 3896
rect 500644 3884 500650 3936
rect 514846 3884 514852 3936
rect 514904 3924 514910 3936
rect 564434 3924 564440 3936
rect 514904 3896 564440 3924
rect 514904 3884 514910 3896
rect 564434 3884 564440 3896
rect 564492 3884 564498 3936
rect 401318 3856 401324 3868
rect 383626 3828 401324 3856
rect 401318 3816 401324 3828
rect 401376 3816 401382 3868
rect 405734 3816 405740 3868
rect 405792 3856 405798 3868
rect 436738 3856 436744 3868
rect 405792 3828 436744 3856
rect 405792 3816 405798 3828
rect 436738 3816 436744 3828
rect 436796 3816 436802 3868
rect 451274 3816 451280 3868
rect 451332 3856 451338 3868
rect 489914 3856 489920 3868
rect 451332 3828 489920 3856
rect 451332 3816 451338 3828
rect 489914 3816 489920 3828
rect 489972 3816 489978 3868
rect 524414 3816 524420 3868
rect 524472 3856 524478 3868
rect 575106 3856 575112 3868
rect 524472 3828 575112 3856
rect 524472 3816 524478 3828
rect 575106 3816 575112 3828
rect 575164 3816 575170 3868
rect 298152 3760 300900 3788
rect 298152 3748 298158 3760
rect 302142 3748 302148 3800
rect 302200 3788 302206 3800
rect 312630 3788 312636 3800
rect 302200 3760 312636 3788
rect 302200 3748 302206 3760
rect 312630 3748 312636 3760
rect 312688 3748 312694 3800
rect 357434 3748 357440 3800
rect 357492 3788 357498 3800
rect 379974 3788 379980 3800
rect 357492 3760 379980 3788
rect 357492 3748 357498 3760
rect 379974 3748 379980 3760
rect 380032 3748 380038 3800
rect 385034 3748 385040 3800
rect 385092 3788 385098 3800
rect 411898 3788 411904 3800
rect 385092 3760 411904 3788
rect 385092 3748 385098 3760
rect 411898 3748 411904 3760
rect 411956 3748 411962 3800
rect 415394 3748 415400 3800
rect 415452 3788 415458 3800
rect 447410 3788 447416 3800
rect 415452 3760 447416 3788
rect 415452 3748 415458 3760
rect 447410 3748 447416 3760
rect 447468 3748 447474 3800
rect 454034 3748 454040 3800
rect 454092 3788 454098 3800
rect 493502 3788 493508 3800
rect 454092 3760 493508 3788
rect 454092 3748 454098 3760
rect 493502 3748 493508 3760
rect 493560 3748 493566 3800
rect 521654 3748 521660 3800
rect 521712 3788 521718 3800
rect 571518 3788 571524 3800
rect 521712 3760 571524 3788
rect 521712 3748 521718 3760
rect 571518 3748 571524 3760
rect 571576 3748 571582 3800
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 49786 3720 49792 3732
rect 20680 3692 49792 3720
rect 20680 3680 20686 3692
rect 49786 3680 49792 3692
rect 49844 3680 49850 3732
rect 53742 3680 53748 3732
rect 53800 3720 53806 3732
rect 78674 3720 78680 3732
rect 53800 3692 78680 3720
rect 53800 3680 53806 3692
rect 78674 3680 78680 3692
rect 78732 3680 78738 3732
rect 84470 3680 84476 3732
rect 84528 3720 84534 3732
rect 101858 3720 101864 3732
rect 84528 3692 101864 3720
rect 84528 3680 84534 3692
rect 101858 3680 101864 3692
rect 101916 3680 101922 3732
rect 110322 3720 110328 3732
rect 104084 3692 110328 3720
rect 8754 3612 8760 3664
rect 8812 3652 8818 3664
rect 40218 3652 40224 3664
rect 8812 3624 40224 3652
rect 8812 3612 8818 3624
rect 40218 3612 40224 3624
rect 40276 3612 40282 3664
rect 43070 3612 43076 3664
rect 43128 3652 43134 3664
rect 69014 3652 69020 3664
rect 43128 3624 69020 3652
rect 43128 3612 43134 3624
rect 69014 3612 69020 3624
rect 69072 3612 69078 3664
rect 71498 3612 71504 3664
rect 71556 3652 71562 3664
rect 93946 3652 93952 3664
rect 71556 3624 93952 3652
rect 71556 3612 71562 3624
rect 93946 3612 93952 3624
rect 94004 3612 94010 3664
rect 96246 3612 96252 3664
rect 96304 3652 96310 3664
rect 103974 3652 103980 3664
rect 96304 3624 103980 3652
rect 96304 3612 96310 3624
rect 103974 3612 103980 3624
rect 104032 3612 104038 3664
rect 13538 3544 13544 3596
rect 13596 3584 13602 3596
rect 44358 3584 44364 3596
rect 13596 3556 44364 3584
rect 13596 3544 13602 3556
rect 44358 3544 44364 3556
rect 44416 3544 44422 3596
rect 46658 3544 46664 3596
rect 46716 3584 46722 3596
rect 71774 3584 71780 3596
rect 46716 3556 71780 3584
rect 46716 3544 46722 3556
rect 71774 3544 71780 3556
rect 71832 3544 71838 3596
rect 73798 3544 73804 3596
rect 73856 3584 73862 3596
rect 95234 3584 95240 3596
rect 73856 3556 95240 3584
rect 73856 3544 73862 3556
rect 95234 3544 95240 3556
rect 95292 3544 95298 3596
rect 104084 3584 104112 3692
rect 110322 3680 110328 3692
rect 110380 3680 110386 3732
rect 114002 3680 114008 3732
rect 114060 3720 114066 3732
rect 129734 3720 129740 3732
rect 114060 3692 129740 3720
rect 114060 3680 114066 3692
rect 129734 3680 129740 3692
rect 129792 3680 129798 3732
rect 130562 3680 130568 3732
rect 130620 3720 130626 3732
rect 137094 3720 137100 3732
rect 130620 3692 137100 3720
rect 130620 3680 130626 3692
rect 137094 3680 137100 3692
rect 137152 3680 137158 3732
rect 140038 3680 140044 3732
rect 140096 3720 140102 3732
rect 146938 3720 146944 3732
rect 140096 3692 146944 3720
rect 140096 3680 140102 3692
rect 146938 3680 146944 3692
rect 146996 3680 147002 3732
rect 149514 3680 149520 3732
rect 149572 3720 149578 3732
rect 157242 3720 157248 3732
rect 149572 3692 157248 3720
rect 149572 3680 149578 3692
rect 157242 3680 157248 3692
rect 157300 3680 157306 3732
rect 157794 3680 157800 3732
rect 157852 3720 157858 3732
rect 165338 3720 165344 3732
rect 157852 3692 165344 3720
rect 157852 3680 157858 3692
rect 165338 3680 165344 3692
rect 165396 3680 165402 3732
rect 189718 3680 189724 3732
rect 189776 3720 189782 3732
rect 194594 3720 194600 3732
rect 189776 3692 194600 3720
rect 189776 3680 189782 3692
rect 194594 3680 194600 3692
rect 194652 3680 194658 3732
rect 199102 3680 199108 3732
rect 199160 3720 199166 3732
rect 202874 3720 202880 3732
rect 199160 3692 202880 3720
rect 199160 3680 199166 3692
rect 202874 3680 202880 3692
rect 202932 3680 202938 3732
rect 286134 3680 286140 3732
rect 286192 3720 286198 3732
rect 294874 3720 294880 3732
rect 286192 3692 294880 3720
rect 286192 3680 286198 3692
rect 294874 3680 294880 3692
rect 294932 3680 294938 3732
rect 295058 3680 295064 3732
rect 295116 3720 295122 3732
rect 304350 3720 304356 3732
rect 295116 3692 304356 3720
rect 295116 3680 295122 3692
rect 304350 3680 304356 3692
rect 304408 3680 304414 3732
rect 305914 3680 305920 3732
rect 305972 3720 305978 3732
rect 317322 3720 317328 3732
rect 305972 3692 317328 3720
rect 305972 3680 305978 3692
rect 317322 3680 317328 3692
rect 317380 3680 317386 3732
rect 358906 3680 358912 3732
rect 358964 3720 358970 3732
rect 382366 3720 382372 3732
rect 358964 3692 382372 3720
rect 358964 3680 358970 3692
rect 382366 3680 382372 3692
rect 382424 3680 382430 3732
rect 397454 3680 397460 3732
rect 397512 3720 397518 3732
rect 426158 3720 426164 3732
rect 397512 3692 426164 3720
rect 397512 3680 397518 3692
rect 426158 3680 426164 3692
rect 426216 3680 426222 3732
rect 427814 3680 427820 3732
rect 427872 3720 427878 3732
rect 461578 3720 461584 3732
rect 427872 3692 461584 3720
rect 427872 3680 427878 3692
rect 461578 3680 461584 3692
rect 461636 3680 461642 3732
rect 463694 3680 463700 3732
rect 463752 3720 463758 3732
rect 504174 3720 504180 3732
rect 463752 3692 504180 3720
rect 463752 3680 463758 3692
rect 504174 3680 504180 3692
rect 504232 3680 504238 3732
rect 529934 3680 529940 3732
rect 529992 3720 529998 3732
rect 580994 3720 581000 3732
rect 529992 3692 581000 3720
rect 529992 3680 529998 3692
rect 580994 3680 581000 3692
rect 581052 3680 581058 3732
rect 106918 3612 106924 3664
rect 106976 3652 106982 3664
rect 124122 3652 124128 3664
rect 106976 3624 124128 3652
rect 106976 3612 106982 3624
rect 124122 3612 124128 3624
rect 124180 3612 124186 3664
rect 154206 3612 154212 3664
rect 154264 3652 154270 3664
rect 160094 3652 160100 3664
rect 154264 3624 160100 3652
rect 154264 3612 154270 3624
rect 160094 3612 160100 3624
rect 160152 3612 160158 3664
rect 170766 3612 170772 3664
rect 170824 3652 170830 3664
rect 177942 3652 177948 3664
rect 170824 3624 177948 3652
rect 170824 3612 170830 3624
rect 177942 3612 177948 3624
rect 178000 3612 178006 3664
rect 253474 3612 253480 3664
rect 253532 3652 253538 3664
rect 255866 3652 255872 3664
rect 253532 3624 255872 3652
rect 253532 3612 253538 3624
rect 255866 3612 255872 3624
rect 255924 3612 255930 3664
rect 259454 3612 259460 3664
rect 259512 3652 259518 3664
rect 264146 3652 264152 3664
rect 259512 3624 264152 3652
rect 259512 3612 259518 3624
rect 264146 3612 264152 3624
rect 264204 3612 264210 3664
rect 267734 3612 267740 3664
rect 267792 3652 267798 3664
rect 273622 3652 273628 3664
rect 267792 3624 273628 3652
rect 267792 3612 267798 3624
rect 273622 3612 273628 3624
rect 273680 3612 273686 3664
rect 278774 3612 278780 3664
rect 278832 3652 278838 3664
rect 286594 3652 286600 3664
rect 278832 3624 286600 3652
rect 278832 3612 278838 3624
rect 286594 3612 286600 3624
rect 286652 3612 286658 3664
rect 288434 3612 288440 3664
rect 288492 3652 288498 3664
rect 298462 3652 298468 3664
rect 288492 3624 298468 3652
rect 288492 3612 288498 3624
rect 298462 3612 298468 3624
rect 298520 3612 298526 3664
rect 303062 3612 303068 3664
rect 303120 3652 303126 3664
rect 313826 3652 313832 3664
rect 303120 3624 313832 3652
rect 303120 3612 303126 3624
rect 313826 3612 313832 3624
rect 313884 3612 313890 3664
rect 345198 3612 345204 3664
rect 345256 3652 345262 3664
rect 346946 3652 346952 3664
rect 345256 3624 346952 3652
rect 345256 3612 345262 3624
rect 346946 3612 346952 3624
rect 347004 3612 347010 3664
rect 363046 3612 363052 3664
rect 363104 3652 363110 3664
rect 387150 3652 387156 3664
rect 363104 3624 387156 3652
rect 363104 3612 363110 3624
rect 387150 3612 387156 3624
rect 387208 3612 387214 3664
rect 393314 3612 393320 3664
rect 393372 3652 393378 3664
rect 422570 3652 422576 3664
rect 393372 3624 422576 3652
rect 393372 3612 393378 3624
rect 422570 3612 422576 3624
rect 422628 3612 422634 3664
rect 434714 3612 434720 3664
rect 434772 3652 434778 3664
rect 471054 3652 471060 3664
rect 434772 3624 471060 3652
rect 434772 3612 434778 3624
rect 471054 3612 471060 3624
rect 471112 3612 471118 3664
rect 476114 3612 476120 3664
rect 476172 3652 476178 3664
rect 518342 3652 518348 3664
rect 476172 3624 518348 3652
rect 476172 3612 476178 3624
rect 518342 3612 518348 3624
rect 518400 3612 518406 3664
rect 527174 3612 527180 3664
rect 527232 3652 527238 3664
rect 578602 3652 578608 3664
rect 527232 3624 578608 3652
rect 527232 3612 527238 3624
rect 578602 3612 578608 3624
rect 578660 3612 578666 3664
rect 99346 3556 104112 3584
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 4798 3516 4804 3528
rect 2924 3488 4804 3516
rect 2924 3476 2930 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 35894 3516 35900 3528
rect 6886 3488 35900 3516
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 6886 3448 6914 3488
rect 35894 3476 35900 3488
rect 35952 3476 35958 3528
rect 35986 3476 35992 3528
rect 36044 3516 36050 3528
rect 63586 3516 63592 3528
rect 36044 3488 63592 3516
rect 36044 3476 36050 3488
rect 63586 3476 63592 3488
rect 63644 3476 63650 3528
rect 70302 3476 70308 3528
rect 70360 3516 70366 3528
rect 92566 3516 92572 3528
rect 70360 3488 92572 3516
rect 70360 3476 70366 3488
rect 92566 3476 92572 3488
rect 92624 3476 92630 3528
rect 4120 3420 6914 3448
rect 4120 3408 4126 3420
rect 38378 3408 38384 3460
rect 38436 3448 38442 3460
rect 64874 3448 64880 3460
rect 38436 3420 64880 3448
rect 38436 3408 38442 3420
rect 64874 3408 64880 3420
rect 64932 3408 64938 3460
rect 66714 3408 66720 3460
rect 66772 3448 66778 3460
rect 89806 3448 89812 3460
rect 66772 3420 89812 3448
rect 66772 3408 66778 3420
rect 89806 3408 89812 3420
rect 89864 3408 89870 3460
rect 91554 3408 91560 3460
rect 91612 3448 91618 3460
rect 99346 3448 99374 3556
rect 104618 3544 104624 3596
rect 104676 3584 104682 3596
rect 121362 3584 121368 3596
rect 104676 3556 121368 3584
rect 104676 3544 104682 3556
rect 121362 3544 121368 3556
rect 121420 3544 121426 3596
rect 156598 3544 156604 3596
rect 156656 3584 156662 3596
rect 162854 3584 162860 3596
rect 156656 3556 162860 3584
rect 156656 3544 156662 3556
rect 162854 3544 162860 3556
rect 162912 3544 162918 3596
rect 180242 3544 180248 3596
rect 180300 3584 180306 3596
rect 186314 3584 186320 3596
rect 180300 3556 186320 3584
rect 180300 3544 180306 3556
rect 186314 3544 186320 3556
rect 186372 3544 186378 3596
rect 234614 3544 234620 3596
rect 234672 3584 234678 3596
rect 235810 3584 235816 3596
rect 234672 3556 235816 3584
rect 234672 3544 234678 3556
rect 235810 3544 235816 3556
rect 235868 3544 235874 3596
rect 258166 3544 258172 3596
rect 258224 3584 258230 3596
rect 262950 3584 262956 3596
rect 258224 3556 262956 3584
rect 258224 3544 258230 3556
rect 262950 3544 262956 3556
rect 263008 3544 263014 3596
rect 266722 3544 266728 3596
rect 266780 3584 266786 3596
rect 272426 3584 272432 3596
rect 266780 3556 272432 3584
rect 266780 3544 266786 3556
rect 272426 3544 272432 3556
rect 272484 3544 272490 3596
rect 285490 3544 285496 3596
rect 285548 3584 285554 3596
rect 292574 3584 292580 3596
rect 285548 3556 292580 3584
rect 285548 3544 285554 3556
rect 292574 3544 292580 3556
rect 292632 3544 292638 3596
rect 293862 3544 293868 3596
rect 293920 3584 293926 3596
rect 303154 3584 303160 3596
rect 293920 3556 303160 3584
rect 293920 3544 293926 3556
rect 303154 3544 303160 3556
rect 303212 3544 303218 3596
rect 304902 3544 304908 3596
rect 304960 3584 304966 3596
rect 315022 3584 315028 3596
rect 304960 3556 315028 3584
rect 304960 3544 304966 3556
rect 315022 3544 315028 3556
rect 315080 3544 315086 3596
rect 331214 3544 331220 3596
rect 331272 3584 331278 3596
rect 333882 3584 333888 3596
rect 331272 3556 333888 3584
rect 331272 3544 331278 3556
rect 333882 3544 333888 3556
rect 333940 3544 333946 3596
rect 334066 3544 334072 3596
rect 334124 3584 334130 3596
rect 344554 3584 344560 3596
rect 334124 3556 344560 3584
rect 334124 3544 334130 3556
rect 344554 3544 344560 3556
rect 344612 3544 344618 3596
rect 346486 3544 346492 3596
rect 346544 3584 346550 3596
rect 348050 3584 348056 3596
rect 346544 3556 348056 3584
rect 346544 3544 346550 3556
rect 348050 3544 348056 3556
rect 348108 3544 348114 3596
rect 349062 3544 349068 3596
rect 349120 3584 349126 3596
rect 351638 3584 351644 3596
rect 349120 3556 351644 3584
rect 349120 3544 349126 3556
rect 351638 3544 351644 3556
rect 351696 3544 351702 3596
rect 353294 3544 353300 3596
rect 353352 3584 353358 3596
rect 355226 3584 355232 3596
rect 353352 3556 355232 3584
rect 353352 3544 353358 3556
rect 355226 3544 355232 3556
rect 355284 3544 355290 3596
rect 362310 3584 362316 3596
rect 355980 3556 362316 3584
rect 101030 3476 101036 3528
rect 101088 3516 101094 3528
rect 118694 3516 118700 3528
rect 101088 3488 118700 3516
rect 101088 3476 101094 3488
rect 118694 3476 118700 3488
rect 118752 3476 118758 3528
rect 119890 3476 119896 3528
rect 119948 3516 119954 3528
rect 135530 3516 135536 3528
rect 119948 3488 135536 3516
rect 119948 3476 119954 3488
rect 135530 3476 135536 3488
rect 135588 3476 135594 3528
rect 142430 3476 142436 3528
rect 142488 3516 142494 3528
rect 149698 3516 149704 3528
rect 142488 3488 149704 3516
rect 142488 3476 142494 3488
rect 149698 3476 149704 3488
rect 149756 3476 149762 3528
rect 153010 3476 153016 3528
rect 153068 3516 153074 3528
rect 158990 3516 158996 3528
rect 153068 3488 158996 3516
rect 153068 3476 153074 3488
rect 158990 3476 158996 3488
rect 159048 3476 159054 3528
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 180702 3516 180708 3528
rect 173216 3488 180708 3516
rect 173216 3476 173222 3488
rect 180702 3476 180708 3488
rect 180760 3476 180766 3528
rect 181438 3476 181444 3528
rect 181496 3516 181502 3528
rect 187694 3516 187700 3528
rect 181496 3488 187700 3516
rect 181496 3476 181502 3488
rect 187694 3476 187700 3488
rect 187752 3476 187758 3528
rect 188522 3476 188528 3528
rect 188580 3516 188586 3528
rect 193214 3516 193220 3528
rect 188580 3488 193220 3516
rect 188580 3476 188586 3488
rect 193214 3476 193220 3488
rect 193272 3476 193278 3528
rect 194410 3476 194416 3528
rect 194468 3516 194474 3528
rect 198734 3516 198740 3528
rect 194468 3488 198740 3516
rect 194468 3476 194474 3488
rect 198734 3476 198740 3488
rect 198792 3476 198798 3528
rect 200298 3476 200304 3528
rect 200356 3516 200362 3528
rect 204346 3516 204352 3528
rect 200356 3488 204352 3516
rect 200356 3476 200362 3488
rect 204346 3476 204352 3488
rect 204404 3476 204410 3528
rect 240226 3476 240232 3528
rect 240284 3516 240290 3528
rect 241698 3516 241704 3528
rect 240284 3488 241704 3516
rect 240284 3476 240290 3488
rect 241698 3476 241704 3488
rect 241756 3476 241762 3528
rect 244642 3476 244648 3528
rect 244700 3516 244706 3528
rect 246390 3516 246396 3528
rect 244700 3488 246396 3516
rect 244700 3476 244706 3488
rect 246390 3476 246396 3488
rect 246448 3476 246454 3528
rect 249794 3476 249800 3528
rect 249852 3516 249858 3528
rect 252370 3516 252376 3528
rect 249852 3488 252376 3516
rect 249852 3476 249858 3488
rect 252370 3476 252376 3488
rect 252428 3476 252434 3528
rect 252462 3476 252468 3528
rect 252520 3516 252526 3528
rect 253474 3516 253480 3528
rect 252520 3488 253480 3516
rect 252520 3476 252526 3488
rect 253474 3476 253480 3488
rect 253532 3476 253538 3528
rect 258074 3476 258080 3528
rect 258132 3516 258138 3528
rect 261754 3516 261760 3528
rect 258132 3488 261760 3516
rect 258132 3476 258138 3488
rect 261754 3476 261760 3488
rect 261812 3476 261818 3528
rect 263502 3476 263508 3528
rect 263560 3516 263566 3528
rect 266538 3516 266544 3528
rect 263560 3488 266544 3516
rect 263560 3476 263566 3488
rect 266538 3476 266544 3488
rect 266596 3476 266602 3528
rect 269114 3476 269120 3528
rect 269172 3516 269178 3528
rect 274818 3516 274824 3528
rect 269172 3488 274824 3516
rect 269172 3476 269178 3488
rect 274818 3476 274824 3488
rect 274876 3476 274882 3528
rect 275830 3476 275836 3528
rect 275888 3516 275894 3528
rect 281902 3516 281908 3528
rect 275888 3488 281908 3516
rect 275888 3476 275894 3488
rect 281902 3476 281908 3488
rect 281960 3476 281966 3528
rect 282730 3476 282736 3528
rect 282788 3516 282794 3528
rect 290182 3516 290188 3528
rect 282788 3488 290188 3516
rect 282788 3476 282794 3488
rect 290182 3476 290188 3488
rect 290240 3476 290246 3528
rect 290826 3476 290832 3528
rect 290884 3516 290890 3528
rect 299658 3516 299664 3528
rect 290884 3488 299664 3516
rect 290884 3476 290890 3488
rect 299658 3476 299664 3488
rect 299716 3476 299722 3528
rect 306374 3476 306380 3528
rect 306432 3516 306438 3528
rect 318518 3516 318524 3528
rect 306432 3488 318524 3516
rect 306432 3476 306438 3488
rect 318518 3476 318524 3488
rect 318576 3476 318582 3528
rect 329650 3476 329656 3528
rect 329708 3516 329714 3528
rect 330386 3516 330392 3528
rect 329708 3488 330392 3516
rect 329708 3476 329714 3488
rect 330386 3476 330392 3488
rect 330444 3476 330450 3528
rect 333238 3476 333244 3528
rect 333296 3516 333302 3528
rect 333296 3488 335354 3516
rect 333296 3476 333302 3488
rect 109678 3448 109684 3460
rect 91612 3420 99374 3448
rect 104176 3420 109684 3448
rect 91612 3408 91618 3420
rect 59630 3340 59636 3392
rect 59688 3380 59694 3392
rect 82814 3380 82820 3392
rect 59688 3352 82820 3380
rect 59688 3340 59694 3352
rect 82814 3340 82820 3352
rect 82872 3340 82878 3392
rect 83274 3340 83280 3392
rect 83332 3380 83338 3392
rect 88886 3380 88892 3392
rect 83332 3352 88892 3380
rect 83332 3340 83338 3352
rect 88886 3340 88892 3352
rect 88944 3340 88950 3392
rect 93946 3340 93952 3392
rect 94004 3380 94010 3392
rect 104176 3380 104204 3420
rect 109678 3408 109684 3420
rect 109736 3408 109742 3460
rect 111610 3408 111616 3460
rect 111668 3448 111674 3460
rect 128262 3448 128268 3460
rect 111668 3420 128268 3448
rect 111668 3408 111674 3420
rect 128262 3408 128268 3420
rect 128320 3408 128326 3460
rect 129366 3408 129372 3460
rect 129424 3448 129430 3460
rect 136542 3448 136548 3460
rect 129424 3420 136548 3448
rect 129424 3408 129430 3420
rect 136542 3408 136548 3420
rect 136600 3408 136606 3460
rect 143534 3408 143540 3460
rect 143592 3448 143598 3460
rect 150434 3448 150440 3460
rect 143592 3420 150440 3448
rect 143592 3408 143598 3420
rect 150434 3408 150440 3420
rect 150492 3408 150498 3460
rect 151814 3408 151820 3460
rect 151872 3448 151878 3460
rect 158806 3448 158812 3460
rect 151872 3420 158812 3448
rect 151872 3408 151878 3420
rect 158806 3408 158812 3420
rect 158864 3408 158870 3460
rect 160094 3408 160100 3460
rect 160152 3448 160158 3460
rect 167270 3448 167276 3460
rect 160152 3420 167276 3448
rect 160152 3408 160158 3420
rect 167270 3408 167276 3420
rect 167328 3408 167334 3460
rect 169570 3408 169576 3460
rect 169628 3448 169634 3460
rect 175274 3448 175280 3460
rect 169628 3420 175280 3448
rect 169628 3408 169634 3420
rect 175274 3408 175280 3420
rect 175332 3408 175338 3460
rect 177850 3408 177856 3460
rect 177908 3448 177914 3460
rect 184842 3448 184848 3460
rect 177908 3420 184848 3448
rect 177908 3408 177914 3420
rect 184842 3408 184848 3420
rect 184900 3408 184906 3460
rect 190822 3408 190828 3460
rect 190880 3448 190886 3460
rect 195974 3448 195980 3460
rect 190880 3420 195980 3448
rect 190880 3408 190886 3420
rect 195974 3408 195980 3420
rect 196032 3408 196038 3460
rect 256602 3408 256608 3460
rect 256660 3448 256666 3460
rect 259454 3448 259460 3460
rect 256660 3420 259460 3448
rect 256660 3408 256666 3420
rect 259454 3408 259460 3420
rect 259512 3408 259518 3460
rect 276750 3408 276756 3460
rect 276808 3448 276814 3460
rect 283098 3448 283104 3460
rect 276808 3420 283104 3448
rect 276808 3408 276814 3420
rect 283098 3408 283104 3420
rect 283156 3408 283162 3460
rect 288526 3408 288532 3460
rect 288584 3448 288590 3460
rect 297266 3448 297272 3460
rect 288584 3420 297272 3448
rect 288584 3408 288590 3420
rect 297266 3408 297272 3420
rect 297324 3408 297330 3460
rect 297450 3408 297456 3460
rect 297508 3448 297514 3460
rect 307938 3448 307944 3460
rect 297508 3420 307944 3448
rect 297508 3408 297514 3420
rect 307938 3408 307944 3420
rect 307996 3408 308002 3460
rect 308030 3408 308036 3460
rect 308088 3448 308094 3460
rect 319714 3448 319720 3460
rect 308088 3420 319720 3448
rect 308088 3408 308094 3420
rect 319714 3408 319720 3420
rect 319772 3408 319778 3460
rect 332686 3408 332692 3460
rect 332744 3448 332750 3460
rect 335078 3448 335084 3460
rect 332744 3420 335084 3448
rect 332744 3408 332750 3420
rect 335078 3408 335084 3420
rect 335136 3408 335142 3460
rect 335326 3448 335354 3488
rect 335538 3476 335544 3528
rect 335596 3516 335602 3528
rect 338666 3516 338672 3528
rect 335596 3488 338672 3516
rect 335596 3476 335602 3488
rect 338666 3476 338672 3488
rect 338724 3476 338730 3528
rect 343726 3476 343732 3528
rect 343784 3516 343790 3528
rect 355980 3516 356008 3556
rect 362310 3544 362316 3556
rect 362368 3544 362374 3596
rect 368382 3544 368388 3596
rect 368440 3584 368446 3596
rect 375190 3584 375196 3596
rect 368440 3556 375196 3584
rect 368440 3544 368446 3556
rect 375190 3544 375196 3556
rect 375248 3544 375254 3596
rect 390646 3584 390652 3596
rect 375392 3556 390652 3584
rect 343784 3488 356008 3516
rect 343784 3476 343790 3488
rect 356054 3476 356060 3528
rect 356112 3516 356118 3528
rect 357526 3516 357532 3528
rect 356112 3488 357532 3516
rect 356112 3476 356118 3488
rect 357526 3476 357532 3488
rect 357584 3476 357590 3528
rect 361758 3476 361764 3528
rect 361816 3516 361822 3528
rect 363506 3516 363512 3528
rect 361816 3488 363512 3516
rect 361816 3476 361822 3488
rect 363506 3476 363512 3488
rect 363564 3476 363570 3528
rect 367186 3476 367192 3528
rect 367244 3516 367250 3528
rect 375392 3516 375420 3556
rect 390646 3544 390652 3556
rect 390704 3544 390710 3596
rect 398834 3544 398840 3596
rect 398892 3584 398898 3596
rect 428458 3584 428464 3596
rect 398892 3556 428464 3584
rect 398892 3544 398898 3556
rect 428458 3544 428464 3556
rect 428516 3544 428522 3596
rect 433334 3544 433340 3596
rect 433392 3584 433398 3596
rect 468662 3584 468668 3596
rect 433392 3556 468668 3584
rect 433392 3544 433398 3556
rect 468662 3544 468668 3556
rect 468720 3544 468726 3596
rect 469214 3544 469220 3596
rect 469272 3584 469278 3596
rect 511258 3584 511264 3596
rect 469272 3556 511264 3584
rect 469272 3544 469278 3556
rect 511258 3544 511264 3556
rect 511316 3544 511322 3596
rect 531406 3544 531412 3596
rect 531464 3584 531470 3596
rect 583386 3584 583392 3596
rect 531464 3556 583392 3584
rect 531464 3544 531470 3556
rect 583386 3544 583392 3556
rect 583444 3544 583450 3596
rect 367244 3488 375420 3516
rect 367244 3476 367250 3488
rect 378134 3476 378140 3528
rect 378192 3516 378198 3528
rect 404814 3516 404820 3528
rect 378192 3488 404820 3516
rect 378192 3476 378198 3488
rect 404814 3476 404820 3488
rect 404872 3476 404878 3528
rect 408494 3476 408500 3528
rect 408552 3516 408558 3528
rect 440326 3516 440332 3528
rect 408552 3488 440332 3516
rect 408552 3476 408558 3488
rect 440326 3476 440332 3488
rect 440384 3476 440390 3528
rect 441614 3476 441620 3528
rect 441672 3516 441678 3528
rect 478138 3516 478144 3528
rect 441672 3488 478144 3516
rect 441672 3476 441678 3488
rect 478138 3476 478144 3488
rect 478196 3476 478202 3528
rect 481634 3476 481640 3528
rect 481692 3516 481698 3528
rect 525426 3516 525432 3528
rect 481692 3488 525432 3516
rect 481692 3476 481698 3488
rect 525426 3476 525432 3488
rect 525484 3476 525490 3528
rect 525794 3476 525800 3528
rect 525852 3516 525858 3528
rect 577406 3516 577412 3528
rect 525852 3488 577412 3516
rect 525852 3476 525858 3488
rect 577406 3476 577412 3488
rect 577464 3476 577470 3528
rect 340966 3448 340972 3460
rect 335326 3420 340972 3448
rect 340966 3408 340972 3420
rect 341024 3408 341030 3460
rect 343634 3408 343640 3460
rect 343692 3448 343698 3460
rect 364610 3448 364616 3460
rect 343692 3420 364616 3448
rect 343692 3408 343698 3420
rect 364610 3408 364616 3420
rect 364668 3408 364674 3460
rect 368290 3408 368296 3460
rect 368348 3448 368354 3460
rect 370590 3448 370596 3460
rect 368348 3420 370596 3448
rect 368348 3408 368354 3420
rect 370590 3408 370596 3420
rect 370648 3408 370654 3460
rect 372614 3408 372620 3460
rect 372672 3448 372678 3460
rect 397730 3448 397736 3460
rect 372672 3420 397736 3448
rect 372672 3408 372678 3420
rect 397730 3408 397736 3420
rect 397788 3408 397794 3460
rect 400214 3408 400220 3460
rect 400272 3448 400278 3460
rect 429654 3448 429660 3460
rect 400272 3420 429660 3448
rect 400272 3408 400278 3420
rect 429654 3408 429660 3420
rect 429712 3408 429718 3460
rect 436094 3408 436100 3460
rect 436152 3448 436158 3460
rect 472250 3448 472256 3460
rect 436152 3420 472256 3448
rect 436152 3408 436158 3420
rect 472250 3408 472256 3420
rect 472308 3408 472314 3460
rect 478966 3408 478972 3460
rect 479024 3448 479030 3460
rect 521838 3448 521844 3460
rect 479024 3420 521844 3448
rect 479024 3408 479030 3420
rect 521838 3408 521844 3420
rect 521896 3408 521902 3460
rect 528554 3408 528560 3460
rect 528612 3448 528618 3460
rect 579798 3448 579804 3460
rect 528612 3420 579804 3448
rect 528612 3408 528618 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 94004 3352 104204 3380
rect 94004 3340 94010 3352
rect 105722 3340 105728 3392
rect 105780 3380 105786 3392
rect 111886 3380 111892 3392
rect 105780 3352 111892 3380
rect 105780 3340 105786 3352
rect 111886 3340 111892 3352
rect 111944 3340 111950 3392
rect 112806 3340 112812 3392
rect 112864 3380 112870 3392
rect 126238 3380 126244 3392
rect 112864 3352 126244 3380
rect 112864 3340 112870 3352
rect 126238 3340 126244 3352
rect 126296 3340 126302 3392
rect 126974 3340 126980 3392
rect 127032 3380 127038 3392
rect 133966 3380 133972 3392
rect 127032 3352 133972 3380
rect 127032 3340 127038 3352
rect 133966 3340 133972 3352
rect 134024 3340 134030 3392
rect 163682 3340 163688 3392
rect 163740 3380 163746 3392
rect 169938 3380 169944 3392
rect 163740 3352 169944 3380
rect 163740 3340 163746 3352
rect 169938 3340 169944 3352
rect 169996 3340 170002 3392
rect 263410 3340 263416 3392
rect 263468 3380 263474 3392
rect 267734 3380 267740 3392
rect 263468 3352 267740 3380
rect 263468 3340 263474 3352
rect 267734 3340 267740 3352
rect 267792 3340 267798 3392
rect 277394 3340 277400 3392
rect 277452 3380 277458 3392
rect 284294 3380 284300 3392
rect 277452 3352 284300 3380
rect 277452 3340 277458 3352
rect 284294 3340 284300 3352
rect 284352 3340 284358 3392
rect 293770 3340 293776 3392
rect 293828 3380 293834 3392
rect 301958 3380 301964 3392
rect 293828 3352 301964 3380
rect 293828 3340 293834 3352
rect 301958 3340 301964 3352
rect 302016 3340 302022 3392
rect 330294 3340 330300 3392
rect 330352 3380 330358 3392
rect 339862 3380 339868 3392
rect 330352 3352 339868 3380
rect 330352 3340 330358 3352
rect 339862 3340 339868 3352
rect 339920 3340 339926 3392
rect 346578 3340 346584 3392
rect 346636 3380 346642 3392
rect 349246 3380 349252 3392
rect 346636 3352 349252 3380
rect 346636 3340 346642 3352
rect 349246 3340 349252 3352
rect 349304 3340 349310 3392
rect 375190 3340 375196 3392
rect 375248 3380 375254 3392
rect 376478 3380 376484 3392
rect 375248 3352 376484 3380
rect 375248 3340 375254 3352
rect 376478 3340 376484 3352
rect 376536 3340 376542 3392
rect 438946 3340 438952 3392
rect 439004 3380 439010 3392
rect 475746 3380 475752 3392
rect 439004 3352 475752 3380
rect 439004 3340 439010 3352
rect 475746 3340 475752 3352
rect 475804 3340 475810 3392
rect 509234 3340 509240 3392
rect 509292 3380 509298 3392
rect 557350 3380 557356 3392
rect 509292 3352 557356 3380
rect 509292 3340 509298 3352
rect 557350 3340 557356 3352
rect 557408 3340 557414 3392
rect 27706 3272 27712 3324
rect 27764 3312 27770 3324
rect 55214 3312 55220 3324
rect 27764 3284 55220 3312
rect 27764 3272 27770 3284
rect 55214 3272 55220 3284
rect 55272 3272 55278 3324
rect 77386 3272 77392 3324
rect 77444 3312 77450 3324
rect 97902 3312 97908 3324
rect 77444 3284 97908 3312
rect 77444 3272 77450 3284
rect 97902 3272 97908 3284
rect 97960 3272 97966 3324
rect 102226 3272 102232 3324
rect 102284 3312 102290 3324
rect 116946 3312 116952 3324
rect 102284 3284 116952 3312
rect 102284 3272 102290 3284
rect 116946 3272 116952 3284
rect 117004 3272 117010 3324
rect 121086 3272 121092 3324
rect 121144 3312 121150 3324
rect 127158 3312 127164 3324
rect 121144 3284 127164 3312
rect 121144 3272 121150 3284
rect 127158 3272 127164 3284
rect 127216 3272 127222 3324
rect 145926 3272 145932 3324
rect 145984 3312 145990 3324
rect 151906 3312 151912 3324
rect 145984 3284 151912 3312
rect 145984 3272 145990 3284
rect 151906 3272 151912 3284
rect 151964 3272 151970 3324
rect 155402 3272 155408 3324
rect 155460 3312 155466 3324
rect 161566 3312 161572 3324
rect 155460 3284 161572 3312
rect 155460 3272 155466 3284
rect 161566 3272 161572 3284
rect 161624 3272 161630 3324
rect 174262 3272 174268 3324
rect 174320 3312 174326 3324
rect 180886 3312 180892 3324
rect 174320 3284 180892 3312
rect 174320 3272 174326 3284
rect 180886 3272 180892 3284
rect 180944 3272 180950 3324
rect 182542 3272 182548 3324
rect 182600 3312 182606 3324
rect 189074 3312 189080 3324
rect 182600 3284 189080 3312
rect 182600 3272 182606 3284
rect 189074 3272 189080 3284
rect 189132 3272 189138 3324
rect 192018 3272 192024 3324
rect 192076 3312 192082 3324
rect 196066 3312 196072 3324
rect 192076 3284 196072 3312
rect 192076 3272 192082 3284
rect 196066 3272 196072 3284
rect 196124 3272 196130 3324
rect 202690 3272 202696 3324
rect 202748 3312 202754 3324
rect 205726 3312 205732 3324
rect 202748 3284 205732 3312
rect 202748 3272 202754 3284
rect 205726 3272 205732 3284
rect 205784 3272 205790 3324
rect 248506 3272 248512 3324
rect 248564 3312 248570 3324
rect 251174 3312 251180 3324
rect 248564 3284 251180 3312
rect 248564 3272 248570 3284
rect 251174 3272 251180 3284
rect 251232 3272 251238 3324
rect 266262 3272 266268 3324
rect 266320 3312 266326 3324
rect 270034 3312 270040 3324
rect 266320 3284 270040 3312
rect 266320 3272 266326 3284
rect 270034 3272 270040 3284
rect 270092 3272 270098 3324
rect 271782 3272 271788 3324
rect 271840 3312 271846 3324
rect 277118 3312 277124 3324
rect 271840 3284 277124 3312
rect 271840 3272 271846 3284
rect 277118 3272 277124 3284
rect 277176 3272 277182 3324
rect 346394 3272 346400 3324
rect 346452 3312 346458 3324
rect 350442 3312 350448 3324
rect 346452 3284 350448 3312
rect 346452 3272 346458 3284
rect 350442 3272 350448 3284
rect 350500 3272 350506 3324
rect 429194 3272 429200 3324
rect 429252 3312 429258 3324
rect 463970 3312 463976 3324
rect 429252 3284 463976 3312
rect 429252 3272 429258 3284
rect 463970 3272 463976 3284
rect 464028 3272 464034 3324
rect 506566 3272 506572 3324
rect 506624 3312 506630 3324
rect 553762 3312 553768 3324
rect 506624 3284 553768 3312
rect 506624 3272 506630 3284
rect 553762 3272 553768 3284
rect 553820 3272 553826 3324
rect 5258 3204 5264 3256
rect 5316 3244 5322 3256
rect 37458 3244 37464 3256
rect 5316 3216 37464 3244
rect 5316 3204 5322 3216
rect 37458 3204 37464 3216
rect 37516 3204 37522 3256
rect 45462 3204 45468 3256
rect 45520 3244 45526 3256
rect 70394 3244 70400 3256
rect 45520 3216 70400 3244
rect 45520 3204 45526 3216
rect 70394 3204 70400 3216
rect 70452 3204 70458 3256
rect 80882 3204 80888 3256
rect 80940 3244 80946 3256
rect 98546 3244 98552 3256
rect 80940 3216 98552 3244
rect 80940 3204 80946 3216
rect 98546 3204 98552 3216
rect 98604 3204 98610 3256
rect 101950 3204 101956 3256
rect 102008 3244 102014 3256
rect 107838 3244 107844 3256
rect 102008 3216 107844 3244
rect 102008 3204 102014 3216
rect 107838 3204 107844 3216
rect 107896 3204 107902 3256
rect 122282 3204 122288 3256
rect 122340 3244 122346 3256
rect 122340 3216 124536 3244
rect 122340 3204 122346 3216
rect 52546 3136 52552 3188
rect 52604 3176 52610 3188
rect 77294 3176 77300 3188
rect 52604 3148 77300 3176
rect 52604 3136 52610 3148
rect 77294 3136 77300 3148
rect 77352 3136 77358 3188
rect 82078 3136 82084 3188
rect 82136 3176 82142 3188
rect 88518 3176 88524 3188
rect 82136 3148 88524 3176
rect 82136 3136 82142 3148
rect 88518 3136 88524 3148
rect 88576 3136 88582 3188
rect 95142 3136 95148 3188
rect 95200 3176 95206 3188
rect 109770 3176 109776 3188
rect 95200 3148 109776 3176
rect 95200 3136 95206 3148
rect 109770 3136 109776 3148
rect 109828 3136 109834 3188
rect 118786 3136 118792 3188
rect 118844 3176 118850 3188
rect 118844 3148 122834 3176
rect 118844 3136 118850 3148
rect 32398 3068 32404 3120
rect 32456 3108 32462 3120
rect 59538 3108 59544 3120
rect 32456 3080 59544 3108
rect 32456 3068 32462 3080
rect 59538 3068 59544 3080
rect 59596 3068 59602 3120
rect 98638 3068 98644 3120
rect 98696 3108 98702 3120
rect 111058 3108 111064 3120
rect 98696 3080 111064 3108
rect 98696 3068 98702 3080
rect 111058 3068 111064 3080
rect 111116 3068 111122 3120
rect 566 3000 572 3052
rect 624 3040 630 3052
rect 2774 3040 2780 3052
rect 624 3012 2780 3040
rect 624 3000 630 3012
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 48958 3000 48964 3052
rect 49016 3040 49022 3052
rect 74718 3040 74724 3052
rect 49016 3012 74724 3040
rect 49016 3000 49022 3012
rect 74718 3000 74724 3012
rect 74776 3000 74782 3052
rect 122806 2972 122834 3148
rect 124508 3108 124536 3216
rect 124674 3204 124680 3256
rect 124732 3244 124738 3256
rect 131114 3244 131120 3256
rect 124732 3216 131120 3244
rect 124732 3204 124738 3216
rect 131114 3204 131120 3216
rect 131172 3204 131178 3256
rect 193214 3204 193220 3256
rect 193272 3244 193278 3256
rect 197354 3244 197360 3256
rect 193272 3216 197360 3244
rect 193272 3204 193278 3216
rect 197354 3204 197360 3216
rect 197412 3204 197418 3256
rect 203886 3204 203892 3256
rect 203944 3244 203950 3256
rect 207106 3244 207112 3256
rect 203944 3216 207112 3244
rect 203944 3204 203950 3216
rect 207106 3204 207112 3216
rect 207164 3204 207170 3256
rect 262122 3204 262128 3256
rect 262180 3244 262186 3256
rect 265342 3244 265348 3256
rect 262180 3216 265348 3244
rect 262180 3204 262186 3216
rect 265342 3204 265348 3216
rect 265400 3204 265406 3256
rect 438854 3204 438860 3256
rect 438912 3244 438918 3256
rect 474550 3244 474556 3256
rect 438912 3216 474556 3244
rect 438912 3204 438918 3216
rect 474550 3204 474556 3216
rect 474608 3204 474614 3256
rect 494054 3204 494060 3256
rect 494112 3244 494118 3256
rect 539594 3244 539600 3256
rect 494112 3216 539600 3244
rect 494112 3204 494118 3216
rect 539594 3204 539600 3216
rect 539652 3204 539658 3256
rect 175458 3136 175464 3188
rect 175516 3176 175522 3188
rect 182174 3176 182180 3188
rect 175516 3148 182180 3176
rect 175516 3136 175522 3148
rect 182174 3136 182180 3148
rect 182232 3136 182238 3188
rect 183738 3136 183744 3188
rect 183796 3176 183802 3188
rect 189166 3176 189172 3188
rect 183796 3148 189172 3176
rect 183796 3136 183802 3148
rect 189166 3136 189172 3148
rect 189224 3136 189230 3188
rect 254762 3136 254768 3188
rect 254820 3176 254826 3188
rect 257062 3176 257068 3188
rect 254820 3148 257068 3176
rect 254820 3136 254826 3148
rect 257062 3136 257068 3148
rect 257120 3136 257126 3188
rect 334158 3136 334164 3188
rect 334216 3176 334222 3188
rect 336274 3176 336280 3188
rect 334216 3148 336280 3176
rect 334216 3136 334222 3148
rect 336274 3136 336280 3148
rect 336332 3136 336338 3188
rect 340782 3136 340788 3188
rect 340840 3176 340846 3188
rect 343358 3176 343364 3188
rect 340840 3148 343364 3176
rect 340840 3136 340846 3148
rect 343358 3136 343364 3148
rect 343416 3136 343422 3188
rect 353386 3136 353392 3188
rect 353444 3176 353450 3188
rect 356330 3176 356336 3188
rect 353444 3148 356336 3176
rect 353444 3136 353450 3148
rect 356330 3136 356336 3148
rect 356388 3136 356394 3188
rect 432046 3136 432052 3188
rect 432104 3176 432110 3188
rect 467466 3176 467472 3188
rect 432104 3148 467472 3176
rect 432104 3136 432110 3148
rect 467466 3136 467472 3148
rect 467524 3136 467530 3188
rect 488534 3136 488540 3188
rect 488592 3176 488598 3188
rect 532510 3176 532516 3188
rect 488592 3148 532516 3176
rect 488592 3136 488598 3148
rect 532510 3136 532516 3148
rect 532568 3136 532574 3188
rect 129642 3108 129648 3120
rect 124508 3080 129648 3108
rect 129642 3068 129648 3080
rect 129700 3068 129706 3120
rect 327074 3068 327080 3120
rect 327132 3108 327138 3120
rect 329190 3108 329196 3120
rect 327132 3080 329196 3108
rect 327132 3068 327138 3080
rect 329190 3068 329196 3080
rect 329248 3068 329254 3120
rect 335446 3068 335452 3120
rect 335504 3108 335510 3120
rect 337470 3108 337476 3120
rect 335504 3080 337476 3108
rect 335504 3068 335510 3080
rect 337470 3068 337476 3080
rect 337528 3068 337534 3120
rect 358630 3068 358636 3120
rect 358688 3108 358694 3120
rect 361114 3108 361120 3120
rect 358688 3080 361120 3108
rect 358688 3068 358694 3080
rect 361114 3068 361120 3080
rect 361172 3068 361178 3120
rect 123478 3000 123484 3052
rect 123536 3040 123542 3052
rect 130378 3040 130384 3052
rect 123536 3012 130384 3040
rect 123536 3000 123542 3012
rect 130378 3000 130384 3012
rect 130436 3000 130442 3052
rect 187326 3000 187332 3052
rect 187384 3040 187390 3052
rect 191926 3040 191932 3052
rect 187384 3012 191932 3040
rect 187384 3000 187390 3012
rect 191926 3000 191932 3012
rect 191984 3000 191990 3052
rect 243262 3000 243268 3052
rect 243320 3040 243326 3052
rect 245194 3040 245200 3052
rect 243320 3012 245200 3040
rect 243320 3000 243326 3012
rect 245194 3000 245200 3012
rect 245252 3000 245258 3052
rect 245838 3000 245844 3052
rect 245896 3040 245902 3052
rect 247586 3040 247592 3052
rect 245896 3012 247592 3040
rect 245896 3000 245902 3012
rect 247586 3000 247592 3012
rect 247644 3000 247650 3052
rect 252278 3000 252284 3052
rect 252336 3040 252342 3052
rect 254670 3040 254676 3052
rect 252336 3012 254676 3040
rect 252336 3000 252342 3012
rect 254670 3000 254676 3012
rect 254728 3000 254734 3052
rect 277670 3000 277676 3052
rect 277728 3040 277734 3052
rect 285398 3040 285404 3052
rect 277728 3012 285404 3040
rect 277728 3000 277734 3012
rect 285398 3000 285404 3012
rect 285456 3000 285462 3052
rect 287330 3000 287336 3052
rect 287388 3040 287394 3052
rect 296070 3040 296076 3052
rect 287388 3012 296076 3040
rect 287388 3000 287394 3012
rect 296070 3000 296076 3012
rect 296128 3000 296134 3052
rect 340414 3000 340420 3052
rect 340472 3040 340478 3052
rect 342162 3040 342168 3052
rect 340472 3012 342168 3040
rect 340472 3000 340478 3012
rect 342162 3000 342168 3012
rect 342220 3000 342226 3052
rect 350534 3000 350540 3052
rect 350592 3040 350598 3052
rect 352834 3040 352840 3052
rect 350592 3012 352840 3040
rect 350592 3000 350598 3012
rect 352834 3000 352840 3012
rect 352892 3000 352898 3052
rect 356238 3000 356244 3052
rect 356296 3040 356302 3052
rect 358722 3040 358728 3052
rect 356296 3012 358728 3040
rect 356296 3000 356302 3012
rect 358722 3000 358728 3012
rect 358780 3000 358786 3052
rect 126882 2972 126888 2984
rect 122806 2944 126888 2972
rect 126882 2932 126888 2944
rect 126940 2932 126946 2984
rect 134150 2932 134156 2984
rect 134208 2972 134214 2984
rect 140866 2972 140872 2984
rect 134208 2944 140872 2972
rect 134208 2932 134214 2944
rect 140866 2932 140872 2944
rect 140924 2932 140930 2984
rect 144730 2932 144736 2984
rect 144788 2972 144794 2984
rect 150710 2972 150716 2984
rect 144788 2944 150716 2972
rect 144788 2932 144794 2944
rect 150710 2932 150716 2944
rect 150768 2932 150774 2984
rect 171962 2932 171968 2984
rect 172020 2972 172026 2984
rect 179322 2972 179328 2984
rect 172020 2944 179328 2972
rect 172020 2932 172026 2944
rect 179322 2932 179328 2944
rect 179380 2932 179386 2984
rect 269206 2932 269212 2984
rect 269264 2972 269270 2984
rect 276014 2972 276020 2984
rect 269264 2944 276020 2972
rect 269264 2932 269270 2944
rect 276014 2932 276020 2944
rect 276072 2932 276078 2984
rect 162486 2864 162492 2916
rect 162544 2904 162550 2916
rect 168466 2904 168472 2916
rect 162544 2876 168472 2904
rect 162544 2864 162550 2876
rect 168466 2864 168472 2876
rect 168524 2864 168530 2916
rect 186130 2864 186136 2916
rect 186188 2904 186194 2916
rect 191834 2904 191840 2916
rect 186188 2876 191840 2904
rect 186188 2864 186194 2876
rect 191834 2864 191840 2876
rect 191892 2864 191898 2916
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 349160 700476 349212 700528
rect 364984 700476 365036 700528
rect 514760 700408 514812 700460
rect 543464 700408 543516 700460
rect 364340 700340 364392 700392
rect 381176 700340 381228 700392
rect 394700 700340 394752 700392
rect 413652 700340 413704 700392
rect 425060 700340 425112 700392
rect 446128 700340 446180 700392
rect 454040 700340 454092 700392
rect 478512 700340 478564 700392
rect 484400 700340 484452 700392
rect 510988 700340 511040 700392
rect 529940 700340 529992 700392
rect 559656 700340 559708 700392
rect 244280 700272 244332 700324
rect 251456 700272 251508 700324
rect 274640 700272 274692 700324
rect 283840 700272 283892 700324
rect 289820 700272 289872 700324
rect 300124 700272 300176 700324
rect 305000 700272 305052 700324
rect 316316 700272 316368 700324
rect 320180 700272 320232 700324
rect 332508 700272 332560 700324
rect 333980 700272 334032 700324
rect 348792 700272 348844 700324
rect 379520 700272 379572 700324
rect 397460 700272 397512 700324
rect 409880 700272 409932 700324
rect 429844 700272 429896 700324
rect 438860 700272 438912 700324
rect 462320 700272 462372 700324
rect 469220 700272 469272 700324
rect 494796 700272 494848 700324
rect 499580 700272 499632 700324
rect 527180 700272 527232 700324
rect 545120 700272 545172 700324
rect 575848 700272 575900 700324
rect 154120 699660 154172 699712
rect 154580 699660 154632 699712
rect 213920 699660 213972 699712
rect 218980 699660 219032 699712
rect 229100 699660 229152 699712
rect 235172 699660 235224 699712
rect 259460 699660 259512 699712
rect 267648 699660 267700 699712
rect 555424 696940 555476 696992
rect 580172 696940 580224 696992
rect 555516 683136 555568 683188
rect 580172 683136 580224 683188
rect 555608 670692 555660 670744
rect 580172 670692 580224 670744
rect 104900 666476 104952 666528
rect 109960 666476 110012 666528
rect 136640 666476 136692 666528
rect 139952 666476 140004 666528
rect 200580 666476 200632 666528
rect 201500 666476 201552 666528
rect 6920 665796 6972 665848
rect 19984 665796 20036 665848
rect 23480 665796 23532 665848
rect 34980 665796 35032 665848
rect 40040 665796 40092 665848
rect 49976 665796 50028 665848
rect 56600 665796 56652 665848
rect 64972 665796 65024 665848
rect 71780 665796 71832 665848
rect 80060 665796 80112 665848
rect 185584 665660 185636 665712
rect 186320 665660 186372 665712
rect 88340 665184 88392 665236
rect 95240 665184 95292 665236
rect 121460 665184 121512 665236
rect 124956 665184 125008 665236
rect 3424 655460 3476 655512
rect 9404 655460 9456 655512
rect 555700 643084 555752 643136
rect 580172 643084 580224 643136
rect 3516 643016 3568 643068
rect 9404 643016 9456 643068
rect 3608 632000 3660 632052
rect 9404 632000 9456 632052
rect 555424 630640 555476 630692
rect 579988 630640 580040 630692
rect 3700 619556 3752 619608
rect 9404 619556 9456 619608
rect 555148 619556 555200 619608
rect 580264 619556 580316 619608
rect 555516 616836 555568 616888
rect 580172 616836 580224 616888
rect 3424 607112 3476 607164
rect 9404 607112 9456 607164
rect 555608 603100 555660 603152
rect 580172 603100 580224 603152
rect 3516 596096 3568 596148
rect 9404 596096 9456 596148
rect 555424 590656 555476 590708
rect 579804 590656 579856 590708
rect 3608 583652 3660 583704
rect 9404 583652 9456 583704
rect 555516 576852 555568 576904
rect 580172 576852 580224 576904
rect 3700 571276 3752 571328
rect 8668 571276 8720 571328
rect 555608 563048 555660 563100
rect 579804 563048 579856 563100
rect 3424 559648 3476 559700
rect 9404 559648 9456 559700
rect 555424 550604 555476 550656
rect 580172 550604 580224 550656
rect 3516 547816 3568 547868
rect 8668 547816 8720 547868
rect 555700 536800 555752 536852
rect 580172 536800 580224 536852
rect 3608 535372 3660 535424
rect 9404 535372 9456 535424
rect 555516 524424 555568 524476
rect 580172 524424 580224 524476
rect 3424 524356 3476 524408
rect 9036 524356 9088 524408
rect 3516 511232 3568 511284
rect 9404 511232 9456 511284
rect 555424 510620 555476 510672
rect 580172 510620 580224 510672
rect 3608 499468 3660 499520
rect 9404 499468 9456 499520
rect 555608 496816 555660 496868
rect 580172 496816 580224 496868
rect 3424 488452 3476 488504
rect 9036 488452 9088 488504
rect 555516 484372 555568 484424
rect 580172 484372 580224 484424
rect 3700 476008 3752 476060
rect 8668 476008 8720 476060
rect 555424 470568 555476 470620
rect 579988 470568 580040 470620
rect 3516 463020 3568 463072
rect 9404 463020 9456 463072
rect 555516 456764 555568 456816
rect 580172 456764 580224 456816
rect 3608 452548 3660 452600
rect 9036 452548 9088 452600
rect 555424 444388 555476 444440
rect 580172 444388 580224 444440
rect 3424 440172 3476 440224
rect 9404 440172 9456 440224
rect 555516 430584 555568 430636
rect 580172 430584 580224 430636
rect 3516 427728 3568 427780
rect 9404 427728 9456 427780
rect 555424 418140 555476 418192
rect 580172 418140 580224 418192
rect 3424 416712 3476 416764
rect 9036 416712 9088 416764
rect 555516 404336 555568 404388
rect 580172 404336 580224 404388
rect 3516 404268 3568 404320
rect 9404 404268 9456 404320
rect 3516 397468 3568 397520
rect 7564 397468 7616 397520
rect 3424 391892 3476 391944
rect 9404 391892 9456 391944
rect 555424 390532 555476 390584
rect 580172 390532 580224 390584
rect 3424 383664 3476 383716
rect 9036 383664 9088 383716
rect 555516 378156 555568 378208
rect 580172 378156 580224 378208
rect 3424 371288 3476 371340
rect 8944 371288 8996 371340
rect 555608 364352 555660 364404
rect 580172 364352 580224 364404
rect 2964 357416 3016 357468
rect 6184 357416 6236 357468
rect 555424 351908 555476 351960
rect 580172 351908 580224 351960
rect 3424 345312 3476 345364
rect 8944 345312 8996 345364
rect 6184 343544 6236 343596
rect 9404 343544 9456 343596
rect 555516 338104 555568 338156
rect 580172 338104 580224 338156
rect 3424 332256 3476 332308
rect 7564 332256 7616 332308
rect 555424 324300 555476 324352
rect 580172 324300 580224 324352
rect 3424 319064 3476 319116
rect 7656 319064 7708 319116
rect 555516 311856 555568 311908
rect 580172 311856 580224 311908
rect 2780 305804 2832 305856
rect 6184 305804 6236 305856
rect 555424 298120 555476 298172
rect 580172 298120 580224 298172
rect 6184 296624 6236 296676
rect 9496 296624 9548 296676
rect 2964 292544 3016 292596
rect 6184 292544 6236 292596
rect 555424 284316 555476 284368
rect 580172 284316 580224 284368
rect 6184 284248 6236 284300
rect 8668 284248 8720 284300
rect 3516 279556 3568 279608
rect 8208 279556 8260 279608
rect 555424 271872 555476 271924
rect 579804 271872 579856 271924
rect 3056 266364 3108 266416
rect 9404 266364 9456 266416
rect 556068 258068 556120 258120
rect 580172 258068 580224 258120
rect 3424 254056 3476 254108
rect 8944 254056 8996 254108
rect 555424 244264 555476 244316
rect 579804 244264 579856 244316
rect 3700 235900 3752 235952
rect 9404 235900 9456 235952
rect 555424 231820 555476 231872
rect 580172 231820 580224 231872
rect 4160 224884 4212 224936
rect 8852 224884 8904 224936
rect 555424 218016 555476 218068
rect 580172 218016 580224 218068
rect 3148 213936 3200 213988
rect 9220 213936 9272 213988
rect 555424 205640 555476 205692
rect 580172 205640 580224 205692
rect 3424 201832 3476 201884
rect 8300 201832 8352 201884
rect 555424 191768 555476 191820
rect 580172 191836 580224 191888
rect 3424 188232 3476 188284
rect 9404 188232 9456 188284
rect 555424 178644 555476 178696
rect 580172 178644 580224 178696
rect 3332 175584 3384 175636
rect 9404 175584 9456 175636
rect 555884 166268 555936 166320
rect 580172 166268 580224 166320
rect 3424 162868 3476 162920
rect 9404 162868 9456 162920
rect 555424 153212 555476 153264
rect 579528 153212 579580 153264
rect 3424 150356 3476 150408
rect 8208 150356 8260 150408
rect 555424 139340 555476 139392
rect 580172 139340 580224 139392
rect 3240 136960 3292 137012
rect 8208 136960 8260 137012
rect 555424 126896 555476 126948
rect 580172 126896 580224 126948
rect 3424 123836 3476 123888
rect 8208 123836 8260 123888
rect 555424 113092 555476 113144
rect 579804 113092 579856 113144
rect 3424 110712 3476 110764
rect 8944 110712 8996 110764
rect 4160 103504 4212 103556
rect 9404 103504 9456 103556
rect 555700 100648 555752 100700
rect 580172 100648 580224 100700
rect 4160 91060 4212 91112
rect 9404 91060 9456 91112
rect 554780 86912 554832 86964
rect 580172 86912 580224 86964
rect 555424 73108 555476 73160
rect 580172 73108 580224 73160
rect 3424 71612 3476 71664
rect 8944 71612 8996 71664
rect 555424 60664 555476 60716
rect 580172 60664 580224 60716
rect 3148 59168 3200 59220
rect 8944 59168 8996 59220
rect 4804 55224 4856 55276
rect 9404 55224 9456 55276
rect 555424 46860 555476 46912
rect 580172 46860 580224 46912
rect 2780 45500 2832 45552
rect 4804 45500 4856 45552
rect 3424 44140 3476 44192
rect 9404 44140 9456 44192
rect 555424 33056 555476 33108
rect 580172 33056 580224 33108
rect 3516 31764 3568 31816
rect 9404 31764 9456 31816
rect 555516 20612 555568 20664
rect 579988 20612 580040 20664
rect 6184 19320 6236 19372
rect 9404 19320 9456 19372
rect 219440 9596 219492 9648
rect 220176 9596 220228 9648
rect 322848 9596 322900 9648
rect 335544 9596 335596 9648
rect 340236 9596 340288 9648
rect 356336 9596 356388 9648
rect 492036 9596 492088 9648
rect 498200 9596 498252 9648
rect 499580 9596 499632 9648
rect 500500 9596 500552 9648
rect 143632 9528 143684 9580
rect 150440 9528 150492 9580
rect 151912 9528 151964 9580
rect 157432 9528 157484 9580
rect 165988 9528 166040 9580
rect 168564 9528 168616 9580
rect 261300 9528 261352 9580
rect 263508 9528 263560 9580
rect 307668 9528 307720 9580
rect 33140 9460 33192 9512
rect 33968 9460 34020 9512
rect 44180 9460 44232 9512
rect 45100 9460 45152 9512
rect 55220 9460 55272 9512
rect 56232 9460 56284 9512
rect 67640 9460 67692 9512
rect 68376 9460 68428 9512
rect 70400 9460 70452 9512
rect 71412 9460 71464 9512
rect 85580 9460 85632 9512
rect 86592 9460 86644 9512
rect 89720 9460 89772 9512
rect 90640 9460 90692 9512
rect 107660 9460 107712 9512
rect 109868 9460 109920 9512
rect 110328 9460 110380 9512
rect 110880 9460 110932 9512
rect 116952 9460 117004 9512
rect 120080 9460 120132 9512
rect 121368 9460 121420 9512
rect 122012 9460 122064 9512
rect 131028 9460 131080 9512
rect 132132 9460 132184 9512
rect 133972 9460 134024 9512
rect 141240 9460 141292 9512
rect 146208 9460 146260 9512
rect 151360 9460 151412 9512
rect 157248 9460 157300 9512
rect 160468 9460 160520 9512
rect 167276 9460 167328 9512
rect 169760 9460 169812 9512
rect 171232 9460 171284 9512
rect 173900 9460 173952 9512
rect 175280 9460 175332 9512
rect 177672 9460 177724 9512
rect 200120 9460 200172 9512
rect 200948 9460 201000 9512
rect 201500 9460 201552 9512
rect 204996 9460 205048 9512
rect 206192 9460 206244 9512
rect 209044 9460 209096 9512
rect 210976 9460 211028 9512
rect 213092 9460 213144 9512
rect 213368 9460 213420 9512
rect 215300 9460 215352 9512
rect 215668 9460 215720 9512
rect 217140 9460 217192 9512
rect 231768 9460 231820 9512
rect 232228 9460 232280 9512
rect 232964 9460 233016 9512
rect 233424 9460 233476 9512
rect 233976 9460 234028 9512
rect 234712 9460 234764 9512
rect 235908 9460 235960 9512
rect 237012 9460 237064 9512
rect 245108 9460 245160 9512
rect 245844 9460 245896 9512
rect 251088 9460 251140 9512
rect 252284 9460 252336 9512
rect 253848 9460 253900 9512
rect 255228 9460 255280 9512
rect 256240 9460 256292 9512
rect 257896 9460 257948 9512
rect 262128 9460 262180 9512
rect 263416 9460 263468 9512
rect 265348 9460 265400 9512
rect 267648 9460 267700 9512
rect 273076 9460 273128 9512
rect 274548 9460 274600 9512
rect 275468 9460 275520 9512
rect 276756 9460 276808 9512
rect 280528 9460 280580 9512
rect 282828 9460 282880 9512
rect 283564 9460 283616 9512
rect 285496 9460 285548 9512
rect 287612 9460 287664 9512
rect 288532 9460 288584 9512
rect 292488 9460 292540 9512
rect 293868 9460 293920 9512
rect 301780 9460 301832 9512
rect 303068 9460 303120 9512
rect 306840 9460 306892 9512
rect 308036 9460 308088 9512
rect 309876 9528 309928 9580
rect 316040 9528 316092 9580
rect 319996 9528 320048 9580
rect 63408 9392 63460 9444
rect 64328 9392 64380 9444
rect 97908 9392 97960 9444
rect 98736 9392 98788 9444
rect 140872 9392 140924 9444
rect 147312 9392 147364 9444
rect 153200 9392 153252 9444
rect 158720 9392 158772 9444
rect 165344 9392 165396 9444
rect 167552 9392 167604 9444
rect 175188 9392 175240 9444
rect 175648 9392 175700 9444
rect 221556 9392 221608 9444
rect 222200 9392 222252 9444
rect 236920 9392 236972 9444
rect 238116 9392 238168 9444
rect 246948 9392 247000 9444
rect 247868 9392 247920 9444
rect 252192 9392 252244 9444
rect 253480 9392 253532 9444
rect 263324 9392 263376 9444
rect 264888 9392 264940 9444
rect 274456 9392 274508 9444
rect 275836 9392 275888 9444
rect 285588 9392 285640 9444
rect 286140 9392 286192 9444
rect 294696 9392 294748 9444
rect 295892 9392 295944 9444
rect 300768 9392 300820 9444
rect 302148 9392 302200 9444
rect 304816 9392 304868 9444
rect 305920 9392 305972 9444
rect 320916 9460 320968 9512
rect 321008 9460 321060 9512
rect 325884 9460 325936 9512
rect 326068 9528 326120 9580
rect 340420 9528 340472 9580
rect 341248 9528 341300 9580
rect 359924 9528 359976 9580
rect 496728 9528 496780 9580
rect 525432 9528 525484 9580
rect 328000 9460 328052 9512
rect 328092 9460 328144 9512
rect 334072 9460 334124 9512
rect 343272 9460 343324 9512
rect 343732 9460 343784 9512
rect 344284 9460 344336 9512
rect 361764 9460 361816 9512
rect 366548 9460 366600 9512
rect 371884 9460 371936 9512
rect 378140 9460 378192 9512
rect 379060 9460 379112 9512
rect 405004 9460 405056 9512
rect 406384 9460 406436 9512
rect 408684 9460 408736 9512
rect 411168 9460 411220 9512
rect 413928 9460 413980 9512
rect 419356 9460 419408 9512
rect 432052 9460 432104 9512
rect 432696 9460 432748 9512
rect 447140 9460 447192 9512
rect 447876 9460 447928 9512
rect 454408 9460 454460 9512
rect 467196 9460 467248 9512
rect 475844 9460 475896 9512
rect 504916 9460 504968 9512
rect 520188 9460 520240 9512
rect 533436 9460 533488 9512
rect 317972 9392 318024 9444
rect 332508 9392 332560 9444
rect 333796 9392 333848 9444
rect 349068 9392 349120 9444
rect 350356 9392 350408 9444
rect 368296 9392 368348 9444
rect 459468 9392 459520 9444
rect 476028 9392 476080 9444
rect 477868 9392 477920 9444
rect 485136 9392 485188 9444
rect 487988 9392 488040 9444
rect 519636 9392 519688 9444
rect 31300 9324 31352 9376
rect 59360 9324 59412 9376
rect 111984 9324 112036 9376
rect 115940 9324 115992 9376
rect 126888 9324 126940 9376
rect 134156 9324 134208 9376
rect 142252 9324 142304 9376
rect 149336 9324 149388 9376
rect 150440 9324 150492 9376
rect 155408 9324 155460 9376
rect 167092 9324 167144 9376
rect 170588 9324 170640 9376
rect 241060 9324 241112 9376
rect 242808 9324 242860 9376
rect 260288 9324 260340 9376
rect 262128 9324 262180 9376
rect 271420 9324 271472 9376
rect 273168 9324 273220 9376
rect 290648 9324 290700 9376
rect 292488 9324 292540 9376
rect 316040 9324 316092 9376
rect 323308 9324 323360 9376
rect 323400 9324 323452 9376
rect 331036 9324 331088 9376
rect 332140 9324 332192 9376
rect 346584 9324 346636 9376
rect 348332 9324 348384 9376
rect 368204 9324 368256 9376
rect 415124 9324 415176 9376
rect 430672 9324 430724 9376
rect 463608 9324 463660 9376
rect 478880 9324 478932 9376
rect 496084 9324 496136 9376
rect 498016 9324 498068 9376
rect 498200 9324 498252 9376
rect 536104 9324 536156 9376
rect 25320 9256 25372 9308
rect 54208 9256 54260 9308
rect 132592 9256 132644 9308
rect 140228 9256 140280 9308
rect 158996 9256 159048 9308
rect 163504 9256 163556 9308
rect 169944 9256 169996 9308
rect 172612 9256 172664 9308
rect 216864 9256 216916 9308
rect 218152 9256 218204 9308
rect 249156 9256 249208 9308
rect 249800 9256 249852 9308
rect 272432 9256 272484 9308
rect 274456 9256 274508 9308
rect 284208 9256 284260 9308
rect 285588 9256 285640 9308
rect 299388 9256 299440 9308
rect 299940 9256 299992 9308
rect 308864 9256 308916 9308
rect 19432 9188 19484 9240
rect 49148 9188 49200 9240
rect 88524 9188 88576 9240
rect 102784 9188 102836 9240
rect 111064 9188 111116 9240
rect 117044 9188 117096 9240
rect 130384 9188 130436 9240
rect 138204 9188 138256 9240
rect 140044 9188 140096 9240
rect 146300 9188 146352 9240
rect 148968 9188 149020 9240
rect 153384 9188 153436 9240
rect 157708 9188 157760 9240
rect 161664 9188 161716 9240
rect 257988 9188 258040 9240
rect 258172 9188 258224 9240
rect 298744 9188 298796 9240
rect 300768 9188 300820 9240
rect 311808 9188 311860 9240
rect 322020 9256 322072 9308
rect 335452 9256 335504 9308
rect 343640 9256 343692 9308
rect 344652 9256 344704 9308
rect 347320 9256 347372 9308
rect 367008 9256 367060 9308
rect 389824 9256 389876 9308
rect 403072 9256 403124 9308
rect 424232 9256 424284 9308
rect 445668 9256 445720 9308
rect 465724 9256 465776 9308
rect 484308 9256 484360 9308
rect 485596 9256 485648 9308
rect 529020 9256 529072 9308
rect 23020 9120 23072 9172
rect 52460 9120 52512 9172
rect 88892 9120 88944 9172
rect 103796 9120 103848 9172
rect 103980 9120 104032 9172
rect 114928 9120 114980 9172
rect 127164 9120 127216 9172
rect 136180 9120 136232 9172
rect 136548 9120 136600 9172
rect 143540 9120 143592 9172
rect 150716 9120 150768 9172
rect 156420 9120 156472 9172
rect 246120 9120 246172 9172
rect 248328 9120 248380 9172
rect 282552 9120 282604 9172
rect 284208 9120 284260 9172
rect 289636 9120 289688 9172
rect 290832 9120 290884 9172
rect 314568 9120 314620 9172
rect 322112 9188 322164 9240
rect 329748 9188 329800 9240
rect 345204 9188 345256 9240
rect 351368 9188 351420 9240
rect 365444 9188 365496 9240
rect 365536 9188 365588 9240
rect 370136 9188 370188 9240
rect 371424 9188 371476 9240
rect 391388 9188 391440 9240
rect 402796 9188 402848 9240
rect 431960 9188 432012 9240
rect 445484 9188 445536 9240
rect 464068 9188 464120 9240
rect 474648 9188 474700 9240
rect 492588 9188 492640 9240
rect 503168 9188 503220 9240
rect 546500 9188 546552 9240
rect 15936 9052 15988 9104
rect 46112 9052 46164 9104
rect 64328 9052 64380 9104
rect 87604 9052 87656 9104
rect 98552 9052 98604 9104
rect 101772 9052 101824 9104
rect 103336 9052 103388 9104
rect 121000 9052 121052 9104
rect 131120 9052 131172 9104
rect 139400 9052 139452 9104
rect 155316 9052 155368 9104
rect 159456 9052 159508 9104
rect 277308 9052 277360 9104
rect 277676 9052 277728 9104
rect 325608 9120 325660 9172
rect 331128 9120 331180 9172
rect 346492 9120 346544 9172
rect 356060 9120 356112 9172
rect 377680 9120 377732 9172
rect 383568 9120 383620 9172
rect 400036 9120 400088 9172
rect 419172 9120 419224 9172
rect 450912 9120 450964 9172
rect 451188 9120 451240 9172
rect 474096 9120 474148 9172
rect 481548 9120 481600 9172
rect 498292 9120 498344 9172
rect 504180 9120 504232 9172
rect 550272 9120 550324 9172
rect 327080 9052 327132 9104
rect 328000 9052 328052 9104
rect 332692 9052 332744 9104
rect 336188 9052 336240 9104
rect 354036 9052 354088 9104
rect 354404 9052 354456 9104
rect 375288 9052 375340 9104
rect 381728 9052 381780 9104
rect 401600 9052 401652 9104
rect 405648 9052 405700 9104
rect 421472 9052 421524 9104
rect 424876 9052 424928 9104
rect 458088 9052 458140 9104
rect 466368 9052 466420 9104
rect 495440 9052 495492 9104
rect 498108 9052 498160 9104
rect 543188 9052 543240 9104
rect 9956 8984 10008 9036
rect 41052 8984 41104 9036
rect 57244 8984 57296 9036
rect 81532 8984 81584 9036
rect 99840 8984 99892 9036
rect 117964 8984 118016 9036
rect 133880 8984 133932 9036
rect 142344 8984 142396 9036
rect 160100 8984 160152 9036
rect 164516 8984 164568 9036
rect 177948 8984 178000 9036
rect 178684 8984 178736 9036
rect 209780 8984 209832 9036
rect 212080 8984 212132 9036
rect 268384 8984 268436 9036
rect 269120 8984 269172 9036
rect 291660 8984 291712 9036
rect 293776 8984 293828 9036
rect 302792 8984 302844 9036
rect 304908 8984 304960 9036
rect 315856 8984 315908 9036
rect 329656 8984 329708 9036
rect 346308 8984 346360 9036
rect 365812 8984 365864 9036
rect 369584 8984 369636 9036
rect 389732 8984 389784 9036
rect 401968 8984 402020 9036
rect 418804 8984 418856 9036
rect 420828 8984 420880 9036
rect 453304 8984 453356 9036
rect 467748 8984 467800 9036
rect 507676 8984 507728 9036
rect 515128 8984 515180 9036
rect 563244 8984 563296 9036
rect 6460 8916 6512 8968
rect 38016 8916 38068 8968
rect 50160 8916 50212 8968
rect 75460 8916 75512 8968
rect 92756 8916 92808 8968
rect 111800 8916 111852 8968
rect 111892 8916 111944 8968
rect 123024 8916 123076 8968
rect 129648 8916 129700 8968
rect 137192 8916 137244 8968
rect 138204 8916 138256 8968
rect 145288 8916 145340 8968
rect 149704 8916 149756 8968
rect 154580 8916 154632 8968
rect 286600 8916 286652 8968
rect 287336 8916 287388 8968
rect 303436 8916 303488 8968
rect 316224 8916 316276 8968
rect 316960 8916 317012 8968
rect 323400 8916 323452 8968
rect 323492 8916 323544 8968
rect 331220 8916 331272 8968
rect 339224 8916 339276 8968
rect 356060 8916 356112 8968
rect 361488 8916 361540 8968
rect 383568 8916 383620 8968
rect 390468 8916 390520 8968
rect 413836 8916 413888 8968
rect 431316 8916 431368 8968
rect 465172 8916 465224 8968
rect 473820 8916 473872 8968
rect 514760 8916 514812 8968
rect 526076 8916 526128 8968
rect 576308 8916 576360 8968
rect 142344 8848 142396 8900
rect 148324 8848 148376 8900
rect 162860 8848 162912 8900
rect 166540 8848 166592 8900
rect 214472 8848 214524 8900
rect 216128 8848 216180 8900
rect 242716 8848 242768 8900
rect 243268 8848 243320 8900
rect 255136 8848 255188 8900
rect 256608 8848 256660 8900
rect 266268 8848 266320 8900
rect 266728 8848 266780 8900
rect 312912 8848 312964 8900
rect 326804 8848 326856 8900
rect 338028 8848 338080 8900
rect 353392 8848 353444 8900
rect 355416 8848 355468 8900
rect 368388 8848 368440 8900
rect 398748 8848 398800 8900
rect 400864 8848 400916 8900
rect 106280 8780 106332 8832
rect 109040 8780 109092 8832
rect 310888 8780 310940 8832
rect 324412 8780 324464 8832
rect 325056 8780 325108 8832
rect 333244 8780 333296 8832
rect 335176 8780 335228 8832
rect 350540 8780 350592 8832
rect 365444 8780 365496 8832
rect 371148 8780 371200 8832
rect 161572 8712 161624 8764
rect 165620 8712 165672 8764
rect 172520 8712 172572 8764
rect 174636 8712 174688 8764
rect 205088 8712 205140 8764
rect 208032 8712 208084 8764
rect 220452 8712 220504 8764
rect 221188 8712 221240 8764
rect 244096 8712 244148 8764
rect 244648 8712 244700 8764
rect 253204 8712 253256 8764
rect 254768 8712 254820 8764
rect 264336 8712 264388 8764
rect 266268 8712 266320 8764
rect 270408 8712 270460 8764
rect 271788 8712 271840 8764
rect 313924 8712 313976 8764
rect 328000 8712 328052 8764
rect 337200 8712 337252 8764
rect 353300 8712 353352 8764
rect 248144 8644 248196 8696
rect 248512 8644 248564 8696
rect 267372 8644 267424 8696
rect 267740 8644 267792 8696
rect 281448 8644 281500 8696
rect 282736 8644 282788 8696
rect 318616 8644 318668 8696
rect 323492 8644 323544 8696
rect 326988 8644 327040 8696
rect 340788 8644 340840 8696
rect 342168 8644 342220 8696
rect 358636 8644 358688 8696
rect 126244 8576 126296 8628
rect 129096 8576 129148 8628
rect 242072 8576 242124 8628
rect 244096 8576 244148 8628
rect 250168 8576 250220 8628
rect 252468 8576 252520 8628
rect 293684 8576 293736 8628
rect 295064 8576 295116 8628
rect 324044 8576 324096 8628
rect 330300 8576 330352 8628
rect 333152 8576 333204 8628
rect 346400 8576 346452 8628
rect 348976 8576 349028 8628
rect 362224 8576 362276 8628
rect 212172 8508 212224 8560
rect 214104 8508 214156 8560
rect 257252 8508 257304 8560
rect 258080 8508 258132 8560
rect 276480 8508 276532 8560
rect 277400 8508 277452 8560
rect 279516 8508 279568 8560
rect 281448 8508 281500 8560
rect 329104 8508 329156 8560
rect 341984 8508 342036 8560
rect 469404 8508 469456 8560
rect 471336 8508 471388 8560
rect 207388 8440 207440 8492
rect 210056 8440 210108 8492
rect 238668 8440 238720 8492
rect 240048 8440 240100 8492
rect 325884 8440 325936 8492
rect 334164 8440 334216 8492
rect 109776 8372 109828 8424
rect 113916 8372 113968 8424
rect 168472 8372 168524 8424
rect 171600 8372 171652 8424
rect 208584 8372 208636 8424
rect 211160 8372 211212 8424
rect 296536 8372 296588 8424
rect 297456 8372 297508 8424
rect 305828 8372 305880 8424
rect 306380 8372 306432 8424
rect 359096 8372 359148 8424
rect 364340 8372 364392 8424
rect 87420 8304 87472 8356
rect 94688 8304 94740 8356
rect 109684 8304 109736 8356
rect 113180 8304 113232 8356
rect 137100 8304 137152 8356
rect 144276 8304 144328 8356
rect 146944 8304 146996 8356
rect 152372 8304 152424 8356
rect 158812 8304 158864 8356
rect 162492 8304 162544 8356
rect 218060 8304 218112 8356
rect 219532 8304 219584 8356
rect 238024 8304 238076 8356
rect 239312 8304 239364 8356
rect 295708 8304 295760 8356
rect 296720 8304 296772 8356
rect 462688 8304 462740 8356
rect 492588 8168 492640 8220
rect 515956 8168 516008 8220
rect 501788 8100 501840 8152
rect 413836 8032 413888 8084
rect 417884 8032 417936 8084
rect 483940 8032 483992 8084
rect 526628 8032 526680 8084
rect 491024 7964 491076 8016
rect 534908 7964 534960 8016
rect 400864 7896 400916 7948
rect 427268 7896 427320 7948
rect 445668 7896 445720 7948
rect 456892 7896 456944 7948
rect 499120 7896 499172 7948
rect 544384 7896 544436 7948
rect 411076 7828 411128 7880
rect 441528 7828 441580 7880
rect 450544 7828 450596 7880
rect 487620 7828 487672 7880
rect 495440 7828 495492 7880
rect 506480 7828 506532 7880
rect 510896 7828 510948 7880
rect 558552 7828 558604 7880
rect 47860 7760 47912 7812
rect 73436 7760 73488 7812
rect 377588 7760 377640 7812
rect 402520 7760 402572 7812
rect 417148 7760 417200 7812
rect 448612 7760 448664 7812
rect 457628 7760 457680 7812
rect 495900 7760 495952 7812
rect 506204 7760 506256 7812
rect 552664 7760 552716 7812
rect 30104 7692 30156 7744
rect 58256 7692 58308 7744
rect 375196 7692 375248 7744
rect 400128 7692 400180 7744
rect 401600 7692 401652 7744
rect 407120 7692 407172 7744
rect 4804 7624 4856 7676
rect 34980 7624 35032 7676
rect 69112 7624 69164 7676
rect 91652 7624 91704 7676
rect 386420 7624 386472 7676
rect 413100 7692 413152 7744
rect 418068 7692 418120 7744
rect 449808 7692 449860 7744
rect 456616 7692 456668 7744
rect 494704 7692 494756 7744
rect 505008 7692 505060 7744
rect 551468 7692 551520 7744
rect 426256 7624 426308 7676
rect 459192 7624 459244 7676
rect 471796 7624 471848 7676
rect 512460 7624 512512 7676
rect 518348 7624 518400 7676
rect 566832 7624 566884 7676
rect 17040 7556 17092 7608
rect 47124 7556 47176 7608
rect 58440 7556 58492 7608
rect 82820 7556 82872 7608
rect 370136 7556 370188 7608
rect 388260 7556 388312 7608
rect 393688 7556 393740 7608
rect 421380 7556 421432 7608
rect 421472 7556 421524 7608
rect 435548 7556 435600 7608
rect 434996 7488 435048 7540
rect 469864 7556 469916 7608
rect 478788 7556 478840 7608
rect 520740 7556 520792 7608
rect 523040 7556 523092 7608
rect 572720 7556 572772 7608
rect 555424 6808 555476 6860
rect 580172 6808 580224 6860
rect 476028 6672 476080 6724
rect 498200 6672 498252 6724
rect 498292 6672 498344 6724
rect 524236 6672 524288 6724
rect 485136 6604 485188 6656
rect 519544 6604 519596 6656
rect 519636 6604 519688 6656
rect 531320 6604 531372 6656
rect 430672 6536 430724 6588
rect 446220 6536 446272 6588
rect 498016 6536 498068 6588
rect 540796 6536 540848 6588
rect 3148 6468 3200 6520
rect 6184 6468 6236 6520
rect 400036 6468 400088 6520
rect 409604 6468 409656 6520
rect 418804 6468 418856 6520
rect 430856 6468 430908 6520
rect 440332 6468 440384 6520
rect 476948 6468 477000 6520
rect 492772 6468 492824 6520
rect 538404 6468 538456 6520
rect 374184 6400 374236 6452
rect 398932 6400 398984 6452
rect 407212 6400 407264 6452
rect 437940 6400 437992 6452
rect 447232 6400 447284 6452
rect 484032 6400 484084 6452
rect 484308 6400 484360 6452
rect 505376 6400 505428 6452
rect 507952 6400 508004 6452
rect 554964 6400 555016 6452
rect 378232 6332 378284 6384
rect 403624 6332 403676 6384
rect 411260 6332 411312 6384
rect 442632 6332 442684 6384
rect 452752 6332 452804 6384
rect 491116 6332 491168 6384
rect 501052 6332 501104 6384
rect 547880 6332 547932 6384
rect 26516 6264 26568 6316
rect 55312 6264 55364 6316
rect 76196 6264 76248 6316
rect 98092 6264 98144 6316
rect 371884 6264 371936 6316
rect 389456 6264 389508 6316
rect 392032 6264 392084 6316
rect 419540 6264 419592 6316
rect 419632 6264 419684 6316
rect 452108 6264 452160 6316
rect 459652 6264 459704 6316
rect 499396 6264 499448 6316
rect 508044 6264 508096 6316
rect 556160 6264 556212 6316
rect 2780 6196 2832 6248
rect 33232 6196 33284 6248
rect 37188 6196 37240 6248
rect 63408 6196 63460 6248
rect 65524 6196 65576 6248
rect 88340 6196 88392 6248
rect 361580 6196 361632 6248
rect 384764 6196 384816 6248
rect 396080 6196 396132 6248
rect 12348 6128 12400 6180
rect 42800 6128 42852 6180
rect 54944 6128 54996 6180
rect 78772 6128 78824 6180
rect 352012 6128 352064 6180
rect 374092 6128 374144 6180
rect 386420 6128 386472 6180
rect 414296 6128 414348 6180
rect 426532 6196 426584 6248
rect 460388 6196 460440 6248
rect 467840 6196 467892 6248
rect 508872 6196 508924 6248
rect 516140 6196 516192 6248
rect 565636 6196 565688 6248
rect 424968 6128 425020 6180
rect 427912 6128 427964 6180
rect 462780 6128 462832 6180
rect 471980 6128 472032 6180
rect 513564 6128 513616 6180
rect 520372 6128 520424 6180
rect 570328 6128 570380 6180
rect 389732 5516 389784 5568
rect 393044 5516 393096 5568
rect 419540 5516 419592 5568
rect 420184 5516 420236 5568
rect 478880 5380 478932 5432
rect 502984 5380 503036 5432
rect 505008 5380 505060 5432
rect 517152 5380 517204 5432
rect 484400 5312 484452 5364
rect 527824 5312 527876 5364
rect 480260 5244 480312 5296
rect 523040 5244 523092 5296
rect 525432 5244 525484 5296
rect 541992 5244 542044 5296
rect 464068 5176 464120 5228
rect 481732 5176 481784 5228
rect 488632 5176 488684 5228
rect 533712 5176 533764 5228
rect 419356 5108 419408 5160
rect 445024 5108 445076 5160
rect 467196 5108 467248 5160
rect 492312 5108 492364 5160
rect 492680 5108 492732 5160
rect 537208 5108 537260 5160
rect 403072 5040 403124 5092
rect 416688 5040 416740 5092
rect 432144 5040 432196 5092
rect 466276 5040 466328 5092
rect 485780 5040 485832 5092
rect 530124 5040 530176 5092
rect 533436 5040 533488 5092
rect 569132 5040 569184 5092
rect 72608 4972 72660 5024
rect 87420 4972 87472 5024
rect 371240 4972 371292 5024
rect 396540 4972 396592 5024
rect 406384 4972 406436 5024
rect 434444 4972 434496 5024
rect 437480 4972 437532 5024
rect 473452 4972 473504 5024
rect 474096 4972 474148 5024
rect 488816 4972 488868 5024
rect 499672 4972 499724 5024
rect 545488 4972 545540 5024
rect 21824 4904 21876 4956
rect 51080 4904 51132 4956
rect 51356 4904 51408 4956
rect 75920 4904 75972 4956
rect 364340 4904 364392 4956
rect 381176 4904 381228 4956
rect 383660 4904 383712 4956
rect 410800 4904 410852 4956
rect 411168 4904 411220 4956
rect 439136 4904 439188 4956
rect 443092 4904 443144 4956
rect 480536 4904 480588 4956
rect 513380 4904 513432 4956
rect 562048 4904 562100 4956
rect 1676 4836 1728 4888
rect 33140 4836 33192 4888
rect 33600 4836 33652 4888
rect 60740 4836 60792 4888
rect 62028 4836 62080 4888
rect 85672 4836 85724 4888
rect 367284 4836 367336 4888
rect 391848 4836 391900 4888
rect 394700 4836 394752 4888
rect 423772 4836 423824 4888
rect 447140 4836 447192 4888
rect 485228 4836 485280 4888
rect 510620 4836 510672 4888
rect 559748 4836 559800 4888
rect 7656 4768 7708 4820
rect 38660 4768 38712 4820
rect 40684 4768 40736 4820
rect 67732 4768 67784 4820
rect 79692 4768 79744 4820
rect 100760 4768 100812 4820
rect 379520 4768 379572 4820
rect 406016 4768 406068 4820
rect 422300 4768 422352 4820
rect 455696 4768 455748 4820
rect 471336 4768 471388 4820
rect 510068 4768 510120 4820
rect 523132 4768 523184 4820
rect 573916 4768 573968 4820
rect 546500 4632 546552 4684
rect 549076 4632 549128 4684
rect 391388 4292 391440 4344
rect 395344 4292 395396 4344
rect 34796 4088 34848 4140
rect 62120 4088 62172 4140
rect 63224 4088 63276 4140
rect 85580 4088 85632 4140
rect 89168 4088 89220 4140
rect 106280 4088 106332 4140
rect 116400 4088 116452 4140
rect 131028 4088 131080 4140
rect 131764 4088 131816 4140
rect 138204 4088 138256 4140
rect 164884 4088 164936 4140
rect 171232 4088 171284 4140
rect 197912 4088 197964 4140
rect 201592 4088 201644 4140
rect 247868 4088 247920 4140
rect 249984 4088 250036 4140
rect 274456 4088 274508 4140
rect 279516 4088 279568 4140
rect 281448 4088 281500 4140
rect 287796 4088 287848 4140
rect 300768 4088 300820 4140
rect 310244 4088 310296 4140
rect 362960 4088 363012 4140
rect 385960 4088 386012 4140
rect 390560 4088 390612 4140
rect 418988 4088 419040 4140
rect 443000 4088 443052 4140
rect 479340 4088 479392 4140
rect 499580 4088 499632 4140
rect 546684 4088 546736 4140
rect 24216 4020 24268 4072
rect 52552 4020 52604 4072
rect 56048 4020 56100 4072
rect 80060 4020 80112 4072
rect 85672 4020 85724 4072
rect 105820 4020 105872 4072
rect 117596 4020 117648 4072
rect 132500 4020 132552 4072
rect 136456 4020 136508 4072
rect 142252 4020 142304 4072
rect 147128 4020 147180 4072
rect 153200 4020 153252 4072
rect 282828 4020 282880 4072
rect 288992 4020 289044 4072
rect 296720 4020 296772 4072
rect 306748 4020 306800 4072
rect 28908 3952 28960 4004
rect 56692 3952 56744 4004
rect 60832 3952 60884 4004
rect 84200 3952 84252 4004
rect 86868 3952 86920 4004
rect 106832 3952 106884 4004
rect 108120 3952 108172 4004
rect 124312 3952 124364 4004
rect 128176 3952 128228 4004
rect 133880 3952 133932 4004
rect 137652 3952 137704 4004
rect 143632 3952 143684 4004
rect 166080 3952 166132 4004
rect 172520 3952 172572 4004
rect 184940 3952 184992 4004
rect 190460 3952 190512 4004
rect 195612 3952 195664 4004
rect 200212 3952 200264 4004
rect 255228 3952 255280 4004
rect 258264 3952 258316 4004
rect 273168 3952 273220 4004
rect 278320 3952 278372 4004
rect 295892 3952 295944 4004
rect 305552 3952 305604 4004
rect 362224 3952 362276 4004
rect 369400 3952 369452 4004
rect 369860 3952 369912 4004
rect 394240 4020 394292 4072
rect 402980 4020 403032 4072
rect 433248 4020 433300 4072
rect 445760 4020 445812 4072
rect 482836 4020 482888 4072
rect 518900 4020 518952 4072
rect 568028 4020 568080 4072
rect 375380 3952 375432 4004
rect 11152 3884 11204 3936
rect 41420 3884 41472 3936
rect 41880 3884 41932 3936
rect 67640 3884 67692 3936
rect 67916 3884 67968 3936
rect 89720 3884 89772 3936
rect 90364 3884 90416 3936
rect 107660 3884 107712 3936
rect 110512 3884 110564 3936
rect 126980 3884 127032 3936
rect 135260 3884 135312 3936
rect 142344 3884 142396 3936
rect 179052 3884 179104 3936
rect 185124 3884 185176 3936
rect 285588 3884 285640 3936
rect 293684 3884 293736 3936
rect 299940 3884 299992 3936
rect 311440 3884 311492 3936
rect 356152 3884 356204 3936
rect 378876 3884 378928 3936
rect 382372 3952 382424 4004
rect 408408 3952 408460 4004
rect 412732 3952 412784 4004
rect 443828 3952 443880 4004
rect 448520 3952 448572 4004
rect 486424 3952 486476 4004
rect 512000 3952 512052 4004
rect 560852 3952 560904 4004
rect 18236 3816 18288 3868
rect 48504 3816 48556 3868
rect 87972 3816 88024 3868
rect 101956 3816 102008 3868
rect 102048 3816 102100 3868
rect 104900 3816 104952 3868
rect 109316 3816 109368 3868
rect 125600 3816 125652 3868
rect 125876 3816 125928 3868
rect 132592 3816 132644 3868
rect 132960 3816 133012 3868
rect 140044 3816 140096 3868
rect 141240 3816 141292 3868
rect 148968 3816 149020 3868
rect 150624 3816 150676 3868
rect 157708 3816 157760 3868
rect 161296 3816 161348 3868
rect 167092 3816 167144 3868
rect 168380 3816 168432 3868
rect 176568 3816 176620 3868
rect 176660 3816 176712 3868
rect 183560 3816 183612 3868
rect 257896 3816 257948 3868
rect 260656 3816 260708 3868
rect 264888 3816 264940 3868
rect 268844 3816 268896 3868
rect 284208 3816 284260 3868
rect 291384 3816 291436 3868
rect 292488 3816 292540 3868
rect 300768 3816 300820 3868
rect 14740 3748 14792 3800
rect 44180 3748 44232 3800
rect 44272 3748 44324 3800
rect 70492 3748 70544 3800
rect 75000 3748 75052 3800
rect 96620 3748 96672 3800
rect 97448 3748 97500 3800
rect 111984 3748 112036 3800
rect 115204 3748 115256 3800
rect 131304 3748 131356 3800
rect 138848 3748 138900 3800
rect 146208 3748 146260 3800
rect 148324 3748 148376 3800
rect 155316 3748 155368 3800
rect 158904 3748 158956 3800
rect 165988 3748 166040 3800
rect 167184 3748 167236 3800
rect 175188 3748 175240 3800
rect 196808 3748 196860 3800
rect 200120 3748 200172 3800
rect 267648 3748 267700 3800
rect 271236 3748 271288 3800
rect 274548 3748 274600 3800
rect 280712 3748 280764 3800
rect 298100 3748 298152 3800
rect 309048 3816 309100 3868
rect 341984 3816 342036 3868
rect 345756 3816 345808 3868
rect 351920 3816 351972 3868
rect 372896 3816 372948 3868
rect 387800 3884 387852 3936
rect 415492 3884 415544 3936
rect 421012 3884 421064 3936
rect 454500 3884 454552 3936
rect 460940 3884 460992 3936
rect 500592 3884 500644 3936
rect 514852 3884 514904 3936
rect 564440 3884 564492 3936
rect 401324 3816 401376 3868
rect 405740 3816 405792 3868
rect 436744 3816 436796 3868
rect 451280 3816 451332 3868
rect 489920 3816 489972 3868
rect 524420 3816 524472 3868
rect 575112 3816 575164 3868
rect 302148 3748 302200 3800
rect 312636 3748 312688 3800
rect 357440 3748 357492 3800
rect 379980 3748 380032 3800
rect 385040 3748 385092 3800
rect 411904 3748 411956 3800
rect 415400 3748 415452 3800
rect 447416 3748 447468 3800
rect 454040 3748 454092 3800
rect 493508 3748 493560 3800
rect 521660 3748 521712 3800
rect 571524 3748 571576 3800
rect 20628 3680 20680 3732
rect 49792 3680 49844 3732
rect 53748 3680 53800 3732
rect 78680 3680 78732 3732
rect 84476 3680 84528 3732
rect 101864 3680 101916 3732
rect 8760 3612 8812 3664
rect 40224 3612 40276 3664
rect 43076 3612 43128 3664
rect 69020 3612 69072 3664
rect 71504 3612 71556 3664
rect 93952 3612 94004 3664
rect 96252 3612 96304 3664
rect 103980 3612 104032 3664
rect 13544 3544 13596 3596
rect 44364 3544 44416 3596
rect 46664 3544 46716 3596
rect 71780 3544 71832 3596
rect 73804 3544 73856 3596
rect 95240 3544 95292 3596
rect 110328 3680 110380 3732
rect 114008 3680 114060 3732
rect 129740 3680 129792 3732
rect 130568 3680 130620 3732
rect 137100 3680 137152 3732
rect 140044 3680 140096 3732
rect 146944 3680 146996 3732
rect 149520 3680 149572 3732
rect 157248 3680 157300 3732
rect 157800 3680 157852 3732
rect 165344 3680 165396 3732
rect 189724 3680 189776 3732
rect 194600 3680 194652 3732
rect 199108 3680 199160 3732
rect 202880 3680 202932 3732
rect 286140 3680 286192 3732
rect 294880 3680 294932 3732
rect 295064 3680 295116 3732
rect 304356 3680 304408 3732
rect 305920 3680 305972 3732
rect 317328 3680 317380 3732
rect 358912 3680 358964 3732
rect 382372 3680 382424 3732
rect 397460 3680 397512 3732
rect 426164 3680 426216 3732
rect 427820 3680 427872 3732
rect 461584 3680 461636 3732
rect 463700 3680 463752 3732
rect 504180 3680 504232 3732
rect 529940 3680 529992 3732
rect 581000 3680 581052 3732
rect 106924 3612 106976 3664
rect 124128 3612 124180 3664
rect 154212 3612 154264 3664
rect 160100 3612 160152 3664
rect 170772 3612 170824 3664
rect 177948 3612 178000 3664
rect 253480 3612 253532 3664
rect 255872 3612 255924 3664
rect 259460 3612 259512 3664
rect 264152 3612 264204 3664
rect 267740 3612 267792 3664
rect 273628 3612 273680 3664
rect 278780 3612 278832 3664
rect 286600 3612 286652 3664
rect 288440 3612 288492 3664
rect 298468 3612 298520 3664
rect 303068 3612 303120 3664
rect 313832 3612 313884 3664
rect 345204 3612 345256 3664
rect 346952 3612 347004 3664
rect 363052 3612 363104 3664
rect 387156 3612 387208 3664
rect 393320 3612 393372 3664
rect 422576 3612 422628 3664
rect 434720 3612 434772 3664
rect 471060 3612 471112 3664
rect 476120 3612 476172 3664
rect 518348 3612 518400 3664
rect 527180 3612 527232 3664
rect 578608 3612 578660 3664
rect 2872 3476 2924 3528
rect 4804 3476 4856 3528
rect 4068 3408 4120 3460
rect 35900 3476 35952 3528
rect 35992 3476 36044 3528
rect 63592 3476 63644 3528
rect 70308 3476 70360 3528
rect 92572 3476 92624 3528
rect 38384 3408 38436 3460
rect 64880 3408 64932 3460
rect 66720 3408 66772 3460
rect 89812 3408 89864 3460
rect 91560 3408 91612 3460
rect 104624 3544 104676 3596
rect 121368 3544 121420 3596
rect 156604 3544 156656 3596
rect 162860 3544 162912 3596
rect 180248 3544 180300 3596
rect 186320 3544 186372 3596
rect 234620 3544 234672 3596
rect 235816 3544 235868 3596
rect 258172 3544 258224 3596
rect 262956 3544 263008 3596
rect 266728 3544 266780 3596
rect 272432 3544 272484 3596
rect 285496 3544 285548 3596
rect 292580 3544 292632 3596
rect 293868 3544 293920 3596
rect 303160 3544 303212 3596
rect 304908 3544 304960 3596
rect 315028 3544 315080 3596
rect 331220 3544 331272 3596
rect 333888 3544 333940 3596
rect 334072 3544 334124 3596
rect 344560 3544 344612 3596
rect 346492 3544 346544 3596
rect 348056 3544 348108 3596
rect 349068 3544 349120 3596
rect 351644 3544 351696 3596
rect 353300 3544 353352 3596
rect 355232 3544 355284 3596
rect 101036 3476 101088 3528
rect 118700 3476 118752 3528
rect 119896 3476 119948 3528
rect 135536 3476 135588 3528
rect 142436 3476 142488 3528
rect 149704 3476 149756 3528
rect 153016 3476 153068 3528
rect 158996 3476 159048 3528
rect 173164 3476 173216 3528
rect 180708 3476 180760 3528
rect 181444 3476 181496 3528
rect 187700 3476 187752 3528
rect 188528 3476 188580 3528
rect 193220 3476 193272 3528
rect 194416 3476 194468 3528
rect 198740 3476 198792 3528
rect 200304 3476 200356 3528
rect 204352 3476 204404 3528
rect 240232 3476 240284 3528
rect 241704 3476 241756 3528
rect 244648 3476 244700 3528
rect 246396 3476 246448 3528
rect 249800 3476 249852 3528
rect 252376 3476 252428 3528
rect 252468 3476 252520 3528
rect 253480 3476 253532 3528
rect 258080 3476 258132 3528
rect 261760 3476 261812 3528
rect 263508 3476 263560 3528
rect 266544 3476 266596 3528
rect 269120 3476 269172 3528
rect 274824 3476 274876 3528
rect 275836 3476 275888 3528
rect 281908 3476 281960 3528
rect 282736 3476 282788 3528
rect 290188 3476 290240 3528
rect 290832 3476 290884 3528
rect 299664 3476 299716 3528
rect 306380 3476 306432 3528
rect 318524 3476 318576 3528
rect 329656 3476 329708 3528
rect 330392 3476 330444 3528
rect 333244 3476 333296 3528
rect 59636 3340 59688 3392
rect 82820 3340 82872 3392
rect 83280 3340 83332 3392
rect 88892 3340 88944 3392
rect 93952 3340 94004 3392
rect 109684 3408 109736 3460
rect 111616 3408 111668 3460
rect 128268 3408 128320 3460
rect 129372 3408 129424 3460
rect 136548 3408 136600 3460
rect 143540 3408 143592 3460
rect 150440 3408 150492 3460
rect 151820 3408 151872 3460
rect 158812 3408 158864 3460
rect 160100 3408 160152 3460
rect 167276 3408 167328 3460
rect 169576 3408 169628 3460
rect 175280 3408 175332 3460
rect 177856 3408 177908 3460
rect 184848 3408 184900 3460
rect 190828 3408 190880 3460
rect 195980 3408 196032 3460
rect 256608 3408 256660 3460
rect 259460 3408 259512 3460
rect 276756 3408 276808 3460
rect 283104 3408 283156 3460
rect 288532 3408 288584 3460
rect 297272 3408 297324 3460
rect 297456 3408 297508 3460
rect 307944 3408 307996 3460
rect 308036 3408 308088 3460
rect 319720 3408 319772 3460
rect 332692 3408 332744 3460
rect 335084 3408 335136 3460
rect 335544 3476 335596 3528
rect 338672 3476 338724 3528
rect 343732 3476 343784 3528
rect 362316 3544 362368 3596
rect 368388 3544 368440 3596
rect 375196 3544 375248 3596
rect 356060 3476 356112 3528
rect 357532 3476 357584 3528
rect 361764 3476 361816 3528
rect 363512 3476 363564 3528
rect 367192 3476 367244 3528
rect 390652 3544 390704 3596
rect 398840 3544 398892 3596
rect 428464 3544 428516 3596
rect 433340 3544 433392 3596
rect 468668 3544 468720 3596
rect 469220 3544 469272 3596
rect 511264 3544 511316 3596
rect 531412 3544 531464 3596
rect 583392 3544 583444 3596
rect 378140 3476 378192 3528
rect 404820 3476 404872 3528
rect 408500 3476 408552 3528
rect 440332 3476 440384 3528
rect 441620 3476 441672 3528
rect 478144 3476 478196 3528
rect 481640 3476 481692 3528
rect 525432 3476 525484 3528
rect 525800 3476 525852 3528
rect 577412 3476 577464 3528
rect 340972 3408 341024 3460
rect 343640 3408 343692 3460
rect 364616 3408 364668 3460
rect 368296 3408 368348 3460
rect 370596 3408 370648 3460
rect 372620 3408 372672 3460
rect 397736 3408 397788 3460
rect 400220 3408 400272 3460
rect 429660 3408 429712 3460
rect 436100 3408 436152 3460
rect 472256 3408 472308 3460
rect 478972 3408 479024 3460
rect 521844 3408 521896 3460
rect 528560 3408 528612 3460
rect 579804 3408 579856 3460
rect 105728 3340 105780 3392
rect 111892 3340 111944 3392
rect 112812 3340 112864 3392
rect 126244 3340 126296 3392
rect 126980 3340 127032 3392
rect 133972 3340 134024 3392
rect 163688 3340 163740 3392
rect 169944 3340 169996 3392
rect 263416 3340 263468 3392
rect 267740 3340 267792 3392
rect 277400 3340 277452 3392
rect 284300 3340 284352 3392
rect 293776 3340 293828 3392
rect 301964 3340 302016 3392
rect 330300 3340 330352 3392
rect 339868 3340 339920 3392
rect 346584 3340 346636 3392
rect 349252 3340 349304 3392
rect 375196 3340 375248 3392
rect 376484 3340 376536 3392
rect 438952 3340 439004 3392
rect 475752 3340 475804 3392
rect 509240 3340 509292 3392
rect 557356 3340 557408 3392
rect 27712 3272 27764 3324
rect 55220 3272 55272 3324
rect 77392 3272 77444 3324
rect 97908 3272 97960 3324
rect 102232 3272 102284 3324
rect 116952 3272 117004 3324
rect 121092 3272 121144 3324
rect 127164 3272 127216 3324
rect 145932 3272 145984 3324
rect 151912 3272 151964 3324
rect 155408 3272 155460 3324
rect 161572 3272 161624 3324
rect 174268 3272 174320 3324
rect 180892 3272 180944 3324
rect 182548 3272 182600 3324
rect 189080 3272 189132 3324
rect 192024 3272 192076 3324
rect 196072 3272 196124 3324
rect 202696 3272 202748 3324
rect 205732 3272 205784 3324
rect 248512 3272 248564 3324
rect 251180 3272 251232 3324
rect 266268 3272 266320 3324
rect 270040 3272 270092 3324
rect 271788 3272 271840 3324
rect 277124 3272 277176 3324
rect 346400 3272 346452 3324
rect 350448 3272 350500 3324
rect 429200 3272 429252 3324
rect 463976 3272 464028 3324
rect 506572 3272 506624 3324
rect 553768 3272 553820 3324
rect 5264 3204 5316 3256
rect 37464 3204 37516 3256
rect 45468 3204 45520 3256
rect 70400 3204 70452 3256
rect 80888 3204 80940 3256
rect 98552 3204 98604 3256
rect 101956 3204 102008 3256
rect 107844 3204 107896 3256
rect 122288 3204 122340 3256
rect 52552 3136 52604 3188
rect 77300 3136 77352 3188
rect 82084 3136 82136 3188
rect 88524 3136 88576 3188
rect 95148 3136 95200 3188
rect 109776 3136 109828 3188
rect 118792 3136 118844 3188
rect 32404 3068 32456 3120
rect 59544 3068 59596 3120
rect 98644 3068 98696 3120
rect 111064 3068 111116 3120
rect 572 3000 624 3052
rect 2780 3000 2832 3052
rect 48964 3000 49016 3052
rect 74724 3000 74776 3052
rect 124680 3204 124732 3256
rect 131120 3204 131172 3256
rect 193220 3204 193272 3256
rect 197360 3204 197412 3256
rect 203892 3204 203944 3256
rect 207112 3204 207164 3256
rect 262128 3204 262180 3256
rect 265348 3204 265400 3256
rect 438860 3204 438912 3256
rect 474556 3204 474608 3256
rect 494060 3204 494112 3256
rect 539600 3204 539652 3256
rect 175464 3136 175516 3188
rect 182180 3136 182232 3188
rect 183744 3136 183796 3188
rect 189172 3136 189224 3188
rect 254768 3136 254820 3188
rect 257068 3136 257120 3188
rect 334164 3136 334216 3188
rect 336280 3136 336332 3188
rect 340788 3136 340840 3188
rect 343364 3136 343416 3188
rect 353392 3136 353444 3188
rect 356336 3136 356388 3188
rect 432052 3136 432104 3188
rect 467472 3136 467524 3188
rect 488540 3136 488592 3188
rect 532516 3136 532568 3188
rect 129648 3068 129700 3120
rect 327080 3068 327132 3120
rect 329196 3068 329248 3120
rect 335452 3068 335504 3120
rect 337476 3068 337528 3120
rect 358636 3068 358688 3120
rect 361120 3068 361172 3120
rect 123484 3000 123536 3052
rect 130384 3000 130436 3052
rect 187332 3000 187384 3052
rect 191932 3000 191984 3052
rect 243268 3000 243320 3052
rect 245200 3000 245252 3052
rect 245844 3000 245896 3052
rect 247592 3000 247644 3052
rect 252284 3000 252336 3052
rect 254676 3000 254728 3052
rect 277676 3000 277728 3052
rect 285404 3000 285456 3052
rect 287336 3000 287388 3052
rect 296076 3000 296128 3052
rect 340420 3000 340472 3052
rect 342168 3000 342220 3052
rect 350540 3000 350592 3052
rect 352840 3000 352892 3052
rect 356244 3000 356296 3052
rect 358728 3000 358780 3052
rect 126888 2932 126940 2984
rect 134156 2932 134208 2984
rect 140872 2932 140924 2984
rect 144736 2932 144788 2984
rect 150716 2932 150768 2984
rect 171968 2932 172020 2984
rect 179328 2932 179380 2984
rect 269212 2932 269264 2984
rect 276020 2932 276072 2984
rect 162492 2864 162544 2916
rect 168472 2864 168524 2916
rect 186136 2864 186188 2916
rect 191840 2864 191892 2916
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 697368 3478 697377
rect 3422 697303 3478 697312
rect 3436 655518 3464 697303
rect 3514 684312 3570 684321
rect 3514 684247 3570 684256
rect 3424 655512 3476 655518
rect 3424 655454 3476 655460
rect 3422 645144 3478 645153
rect 3422 645079 3478 645088
rect 3436 607170 3464 645079
rect 3528 643074 3556 684247
rect 3606 671256 3662 671265
rect 3606 671191 3662 671200
rect 3516 643068 3568 643074
rect 3516 643010 3568 643016
rect 3514 632088 3570 632097
rect 3620 632058 3648 671191
rect 6932 665854 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 23492 665854 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 40052 665854 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 56796 683114 56824 703520
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 56612 683086 56824 683114
rect 56612 665854 56640 683086
rect 71792 665854 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 6920 665848 6972 665854
rect 6920 665790 6972 665796
rect 19984 665848 20036 665854
rect 19984 665790 20036 665796
rect 23480 665848 23532 665854
rect 23480 665790 23532 665796
rect 34980 665848 35032 665854
rect 34980 665790 35032 665796
rect 40040 665848 40092 665854
rect 40040 665790 40092 665796
rect 49976 665848 50028 665854
rect 49976 665790 50028 665796
rect 56600 665848 56652 665854
rect 56600 665790 56652 665796
rect 64972 665848 65024 665854
rect 64972 665790 65024 665796
rect 71780 665848 71832 665854
rect 71780 665790 71832 665796
rect 80060 665848 80112 665854
rect 80060 665790 80112 665796
rect 19996 663490 20024 665790
rect 34992 663490 35020 665790
rect 49988 663490 50016 665790
rect 64984 663490 65012 665790
rect 80072 663490 80100 665790
rect 88352 665242 88380 702406
rect 104912 666534 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 121656 683114 121684 703520
rect 121472 683086 121684 683114
rect 104900 666528 104952 666534
rect 104900 666470 104952 666476
rect 109960 666528 110012 666534
rect 109960 666470 110012 666476
rect 88340 665236 88392 665242
rect 88340 665178 88392 665184
rect 95240 665236 95292 665242
rect 95240 665178 95292 665184
rect 95252 663490 95280 665178
rect 109972 663490 110000 666470
rect 121472 665242 121500 683086
rect 136652 666534 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 699718 154160 703520
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 154120 699712 154172 699718
rect 154120 699654 154172 699660
rect 154580 699712 154632 699718
rect 154580 699654 154632 699660
rect 154592 673454 154620 699654
rect 169772 673454 169800 702406
rect 186516 683114 186544 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 186332 683086 186544 683114
rect 154592 673426 154896 673454
rect 169772 673426 169892 673454
rect 136640 666528 136692 666534
rect 136640 666470 136692 666476
rect 139952 666528 140004 666534
rect 139952 666470 140004 666476
rect 121460 665236 121512 665242
rect 121460 665178 121512 665184
rect 124956 665236 125008 665242
rect 124956 665178 125008 665184
rect 124968 663490 124996 665178
rect 139964 663490 139992 666470
rect 154868 663490 154896 673426
rect 169864 663490 169892 673426
rect 186332 665718 186360 683086
rect 201512 666534 201540 702986
rect 218992 699718 219020 703520
rect 235184 699718 235212 703520
rect 251468 700330 251496 703520
rect 244280 700324 244332 700330
rect 244280 700266 244332 700272
rect 251456 700324 251508 700330
rect 251456 700266 251508 700272
rect 213920 699712 213972 699718
rect 213920 699654 213972 699660
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 229100 699712 229152 699718
rect 229100 699654 229152 699660
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 213932 673454 213960 699654
rect 229112 673454 229140 699654
rect 244292 673454 244320 700266
rect 267660 699718 267688 703520
rect 283852 700330 283880 703520
rect 300136 700330 300164 703520
rect 316328 700330 316356 703520
rect 332520 700330 332548 703520
rect 348804 700330 348832 703520
rect 364996 700534 365024 703520
rect 349160 700528 349212 700534
rect 349160 700470 349212 700476
rect 364984 700528 365036 700534
rect 364984 700470 365036 700476
rect 274640 700324 274692 700330
rect 274640 700266 274692 700272
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 289820 700324 289872 700330
rect 289820 700266 289872 700272
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 305000 700324 305052 700330
rect 305000 700266 305052 700272
rect 316316 700324 316368 700330
rect 316316 700266 316368 700272
rect 320180 700324 320232 700330
rect 320180 700266 320232 700272
rect 332508 700324 332560 700330
rect 332508 700266 332560 700272
rect 333980 700324 334032 700330
rect 333980 700266 334032 700272
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 259460 699712 259512 699718
rect 259460 699654 259512 699660
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 259472 673454 259500 699654
rect 274652 673454 274680 700266
rect 213932 673426 214880 673454
rect 229112 673426 229876 673454
rect 244292 673426 244872 673454
rect 259472 673426 259868 673454
rect 274652 673426 274864 673454
rect 200580 666528 200632 666534
rect 200580 666470 200632 666476
rect 201500 666528 201552 666534
rect 201500 666470 201552 666476
rect 185584 665712 185636 665718
rect 185584 665654 185636 665660
rect 186320 665712 186372 665718
rect 186320 665654 186372 665660
rect 185596 663490 185624 665654
rect 200592 663490 200620 666470
rect 19996 663462 20332 663490
rect 34992 663462 35328 663490
rect 49988 663462 50324 663490
rect 64984 663462 65320 663490
rect 80072 663462 80316 663490
rect 95252 663462 95312 663490
rect 109972 663462 110308 663490
rect 124968 663462 125304 663490
rect 139964 663462 140300 663490
rect 154868 663462 155296 663490
rect 169864 663462 170292 663490
rect 185288 663462 185624 663490
rect 200284 663462 200620 663490
rect 214852 663490 214880 673426
rect 229848 663490 229876 673426
rect 244844 663490 244872 673426
rect 259840 663490 259868 673426
rect 274836 663490 274864 673426
rect 289832 663490 289860 700266
rect 305012 663490 305040 700266
rect 320192 663490 320220 700266
rect 333992 673454 334020 700266
rect 349172 673454 349200 700470
rect 381188 700398 381216 703520
rect 364340 700392 364392 700398
rect 364340 700334 364392 700340
rect 381176 700392 381228 700398
rect 381176 700334 381228 700340
rect 394700 700392 394752 700398
rect 394700 700334 394752 700340
rect 364352 673454 364380 700334
rect 379520 700324 379572 700330
rect 379520 700266 379572 700272
rect 379532 673454 379560 700266
rect 394712 673454 394740 700334
rect 397472 700330 397500 703520
rect 413664 700398 413692 703520
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 425060 700392 425112 700398
rect 425060 700334 425112 700340
rect 397460 700324 397512 700330
rect 397460 700266 397512 700272
rect 409880 700324 409932 700330
rect 409880 700266 409932 700272
rect 333992 673426 334848 673454
rect 349172 673426 349844 673454
rect 364352 673426 364840 673454
rect 379532 673426 379836 673454
rect 394712 673426 394832 673454
rect 334820 663490 334848 673426
rect 349816 663490 349844 673426
rect 364812 663490 364840 673426
rect 379808 663490 379836 673426
rect 394804 663490 394832 673426
rect 409892 663490 409920 700266
rect 425072 663490 425100 700334
rect 429856 700330 429884 703520
rect 446140 700398 446168 703520
rect 446128 700392 446180 700398
rect 446128 700334 446180 700340
rect 454040 700392 454092 700398
rect 454040 700334 454092 700340
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 438860 700324 438912 700330
rect 438860 700266 438912 700272
rect 438872 673454 438900 700266
rect 454052 673454 454080 700334
rect 462332 700330 462360 703520
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 484400 700392 484452 700398
rect 484400 700334 484452 700340
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 469220 700324 469272 700330
rect 469220 700266 469272 700272
rect 469232 673454 469260 700266
rect 484412 673454 484440 700334
rect 494808 700330 494836 703520
rect 511000 700398 511028 703520
rect 514760 700460 514812 700466
rect 514760 700402 514812 700408
rect 510988 700392 511040 700398
rect 510988 700334 511040 700340
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 499580 700324 499632 700330
rect 499580 700266 499632 700272
rect 499592 673454 499620 700266
rect 438872 673426 439820 673454
rect 454052 673426 454816 673454
rect 469232 673426 469812 673454
rect 484412 673426 484808 673454
rect 499592 673426 499804 673454
rect 439792 663490 439820 673426
rect 454788 663490 454816 673426
rect 469784 663490 469812 673426
rect 484780 663490 484808 673426
rect 499776 663490 499804 673426
rect 514772 663490 514800 700402
rect 527192 700330 527220 703520
rect 543476 700466 543504 703520
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 559668 700398 559696 703520
rect 529940 700392 529992 700398
rect 529940 700334 529992 700340
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 529952 663490 529980 700334
rect 575860 700330 575888 703520
rect 545120 700324 545172 700330
rect 545120 700266 545172 700272
rect 575848 700324 575900 700330
rect 575848 700266 575900 700272
rect 545132 663490 545160 700266
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 555424 696992 555476 696998
rect 555424 696934 555476 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 214852 663462 215280 663490
rect 229848 663462 230276 663490
rect 244844 663462 245272 663490
rect 259840 663462 260268 663490
rect 274836 663462 275264 663490
rect 289832 663462 290260 663490
rect 305012 663462 305256 663490
rect 320192 663462 320252 663490
rect 334820 663462 335248 663490
rect 349816 663462 350244 663490
rect 364812 663462 365240 663490
rect 379808 663462 380236 663490
rect 394804 663462 395232 663490
rect 409892 663462 410228 663490
rect 425072 663462 425224 663490
rect 439792 663462 440220 663490
rect 454788 663462 455216 663490
rect 469784 663462 470212 663490
rect 484780 663462 485208 663490
rect 499776 663462 500204 663490
rect 514772 663462 515200 663490
rect 529952 663462 530196 663490
rect 545132 663462 545192 663490
rect 3698 658200 3754 658209
rect 3698 658135 3754 658144
rect 3514 632023 3570 632032
rect 3608 632052 3660 632058
rect 3424 607164 3476 607170
rect 3424 607106 3476 607112
rect 3528 596154 3556 632023
rect 3608 631994 3660 632000
rect 3712 619614 3740 658135
rect 555436 655897 555464 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 555516 683188 555568 683194
rect 555516 683130 555568 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 555422 655888 555478 655897
rect 555422 655823 555478 655832
rect 9404 655512 9456 655518
rect 9404 655454 9456 655460
rect 9416 654809 9444 655454
rect 9402 654800 9458 654809
rect 9402 654735 9458 654744
rect 555528 643657 555556 683130
rect 555608 670744 555660 670750
rect 580172 670744 580224 670750
rect 555608 670686 555660 670692
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 555514 643648 555570 643657
rect 555514 643583 555570 643592
rect 9404 643068 9456 643074
rect 9404 643010 9456 643016
rect 9416 642841 9444 643010
rect 9402 642832 9458 642841
rect 9402 642767 9458 642776
rect 9404 632052 9456 632058
rect 9404 631994 9456 632000
rect 9416 630873 9444 631994
rect 555620 631417 555648 670686
rect 580170 670647 580226 670656
rect 580262 657384 580318 657393
rect 580262 657319 580318 657328
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 555700 643136 555752 643142
rect 555700 643078 555752 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 555606 631408 555662 631417
rect 555606 631343 555662 631352
rect 9402 630864 9458 630873
rect 9402 630799 9458 630808
rect 555424 630692 555476 630698
rect 555424 630634 555476 630640
rect 3700 619608 3752 619614
rect 3700 619550 3752 619556
rect 9404 619608 9456 619614
rect 9404 619550 9456 619556
rect 555148 619608 555200 619614
rect 555148 619550 555200 619556
rect 3606 619168 3662 619177
rect 3606 619103 3662 619112
rect 3516 596148 3568 596154
rect 3516 596090 3568 596096
rect 3422 593056 3478 593065
rect 3422 592991 3478 593000
rect 3436 559706 3464 592991
rect 3620 583710 3648 619103
rect 9416 618905 9444 619550
rect 555160 619177 555188 619550
rect 555146 619168 555202 619177
rect 555146 619103 555202 619112
rect 9402 618896 9458 618905
rect 9402 618831 9458 618840
rect 9404 607164 9456 607170
rect 9404 607106 9456 607112
rect 9416 606937 9444 607106
rect 9402 606928 9458 606937
rect 9402 606863 9458 606872
rect 3698 606112 3754 606121
rect 3698 606047 3754 606056
rect 3608 583704 3660 583710
rect 3608 583646 3660 583652
rect 3514 580000 3570 580009
rect 3514 579935 3570 579944
rect 3424 559700 3476 559706
rect 3424 559642 3476 559648
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 524414 3464 553823
rect 3528 547874 3556 579935
rect 3712 571334 3740 606047
rect 9404 596148 9456 596154
rect 9404 596090 9456 596096
rect 9416 594969 9444 596090
rect 9402 594960 9458 594969
rect 9402 594895 9458 594904
rect 555436 594697 555464 630634
rect 555516 616888 555568 616894
rect 555516 616830 555568 616836
rect 555422 594688 555478 594697
rect 555422 594623 555478 594632
rect 555424 590708 555476 590714
rect 555424 590650 555476 590656
rect 9404 583704 9456 583710
rect 9404 583646 9456 583652
rect 9416 583001 9444 583646
rect 9402 582992 9458 583001
rect 9402 582927 9458 582936
rect 3700 571328 3752 571334
rect 3700 571270 3752 571276
rect 8668 571328 8720 571334
rect 8668 571270 8720 571276
rect 8680 571033 8708 571270
rect 8666 571024 8722 571033
rect 8666 570959 8722 570968
rect 3606 566944 3662 566953
rect 3606 566879 3662 566888
rect 3516 547868 3568 547874
rect 3516 547810 3568 547816
rect 3514 540832 3570 540841
rect 3514 540767 3570 540776
rect 3424 524408 3476 524414
rect 3424 524350 3476 524356
rect 3422 514856 3478 514865
rect 3422 514791 3478 514800
rect 3436 488510 3464 514791
rect 3528 511290 3556 540767
rect 3620 535430 3648 566879
rect 9404 559700 9456 559706
rect 9404 559642 9456 559648
rect 9416 559065 9444 559642
rect 9402 559056 9458 559065
rect 9402 558991 9458 559000
rect 555436 557977 555464 590650
rect 555528 582457 555556 616830
rect 555712 606937 555740 643078
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580276 619614 580304 657319
rect 580264 619608 580316 619614
rect 580264 619550 580316 619556
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 555698 606928 555754 606937
rect 555698 606863 555754 606872
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 555608 603152 555660 603158
rect 555608 603094 555660 603100
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 555514 582448 555570 582457
rect 555514 582383 555570 582392
rect 555516 576904 555568 576910
rect 555516 576846 555568 576852
rect 555422 557968 555478 557977
rect 555422 557903 555478 557912
rect 555424 550656 555476 550662
rect 555424 550598 555476 550604
rect 8668 547868 8720 547874
rect 8668 547810 8720 547816
rect 8680 547097 8708 547810
rect 8666 547088 8722 547097
rect 8666 547023 8722 547032
rect 3608 535424 3660 535430
rect 3608 535366 3660 535372
rect 9404 535424 9456 535430
rect 9404 535366 9456 535372
rect 9416 535129 9444 535366
rect 9402 535120 9458 535129
rect 9402 535055 9458 535064
rect 3606 527912 3662 527921
rect 3606 527847 3662 527856
rect 3516 511284 3568 511290
rect 3516 511226 3568 511232
rect 3620 499526 3648 527847
rect 9036 524408 9088 524414
rect 9036 524350 9088 524356
rect 9048 523161 9076 524350
rect 9034 523152 9090 523161
rect 9034 523087 9090 523096
rect 555436 521257 555464 550598
rect 555528 545737 555556 576846
rect 555620 570217 555648 603094
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 555606 570208 555662 570217
rect 555606 570143 555662 570152
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 555608 563100 555660 563106
rect 555608 563042 555660 563048
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 555514 545728 555570 545737
rect 555514 545663 555570 545672
rect 555620 533497 555648 563042
rect 580170 551168 580226 551177
rect 580170 551103 580226 551112
rect 580184 550662 580212 551103
rect 580172 550656 580224 550662
rect 580172 550598 580224 550604
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 555700 536852 555752 536858
rect 555700 536794 555752 536800
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 555606 533488 555662 533497
rect 555606 533423 555662 533432
rect 555516 524476 555568 524482
rect 555516 524418 555568 524424
rect 555422 521248 555478 521257
rect 555422 521183 555478 521192
rect 9404 511284 9456 511290
rect 9404 511226 9456 511232
rect 9416 511193 9444 511226
rect 9402 511184 9458 511193
rect 9402 511119 9458 511128
rect 555424 510672 555476 510678
rect 555424 510614 555476 510620
rect 3698 501800 3754 501809
rect 3698 501735 3754 501744
rect 3608 499520 3660 499526
rect 3608 499462 3660 499468
rect 3514 488744 3570 488753
rect 3514 488679 3570 488688
rect 3424 488504 3476 488510
rect 3424 488446 3476 488452
rect 3528 463078 3556 488679
rect 3712 476066 3740 501735
rect 9404 499520 9456 499526
rect 9404 499462 9456 499468
rect 9416 499225 9444 499462
rect 9402 499216 9458 499225
rect 9402 499151 9458 499160
rect 9036 488504 9088 488510
rect 9036 488446 9088 488452
rect 9048 487257 9076 488446
rect 9034 487248 9090 487257
rect 9034 487183 9090 487192
rect 555436 484537 555464 510614
rect 555528 496777 555556 524418
rect 555712 509017 555740 536794
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 555698 509008 555754 509017
rect 555698 508943 555754 508952
rect 580170 497992 580226 498001
rect 580170 497927 580226 497936
rect 580184 496874 580212 497927
rect 555608 496868 555660 496874
rect 555608 496810 555660 496816
rect 580172 496868 580224 496874
rect 580172 496810 580224 496816
rect 555514 496768 555570 496777
rect 555514 496703 555570 496712
rect 555422 484528 555478 484537
rect 555422 484463 555478 484472
rect 555516 484424 555568 484430
rect 555516 484366 555568 484372
rect 3700 476060 3752 476066
rect 3700 476002 3752 476008
rect 8668 476060 8720 476066
rect 8668 476002 8720 476008
rect 3606 475688 3662 475697
rect 3606 475623 3662 475632
rect 3516 463072 3568 463078
rect 3516 463014 3568 463020
rect 3422 462632 3478 462641
rect 3422 462567 3478 462576
rect 3436 440230 3464 462567
rect 3620 452606 3648 475623
rect 8680 475289 8708 476002
rect 8666 475280 8722 475289
rect 8666 475215 8722 475224
rect 555424 470620 555476 470626
rect 555424 470562 555476 470568
rect 9402 463312 9458 463321
rect 9402 463247 9458 463256
rect 9416 463078 9444 463247
rect 9404 463072 9456 463078
rect 9404 463014 9456 463020
rect 3608 452600 3660 452606
rect 3608 452542 3660 452548
rect 9036 452600 9088 452606
rect 9036 452542 9088 452548
rect 9048 451353 9076 452542
rect 9034 451344 9090 451353
rect 9034 451279 9090 451288
rect 3514 449576 3570 449585
rect 3514 449511 3570 449520
rect 3424 440224 3476 440230
rect 3424 440166 3476 440172
rect 3422 436656 3478 436665
rect 3422 436591 3478 436600
rect 3436 416770 3464 436591
rect 3528 427786 3556 449511
rect 555436 447817 555464 470562
rect 555528 460057 555556 484366
rect 555620 472297 555648 496810
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 555606 472288 555662 472297
rect 555606 472223 555662 472232
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 555514 460048 555570 460057
rect 555514 459983 555570 459992
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 555516 456816 555568 456822
rect 555516 456758 555568 456764
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 555422 447808 555478 447817
rect 555422 447743 555478 447752
rect 555424 444440 555476 444446
rect 555424 444382 555476 444388
rect 9404 440224 9456 440230
rect 9404 440166 9456 440172
rect 9416 439385 9444 440166
rect 9402 439376 9458 439385
rect 9402 439311 9458 439320
rect 3516 427780 3568 427786
rect 3516 427722 3568 427728
rect 9404 427780 9456 427786
rect 9404 427722 9456 427728
rect 9416 427417 9444 427722
rect 9402 427408 9458 427417
rect 9402 427343 9458 427352
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3424 416764 3476 416770
rect 3424 416706 3476 416712
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3436 391950 3464 410479
rect 3528 404326 3556 423535
rect 555436 423337 555464 444382
rect 555528 435577 555556 456758
rect 580170 444816 580226 444825
rect 580170 444751 580226 444760
rect 580184 444446 580212 444751
rect 580172 444440 580224 444446
rect 580172 444382 580224 444388
rect 555514 435568 555570 435577
rect 555514 435503 555570 435512
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 555516 430636 555568 430642
rect 555516 430578 555568 430584
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 555422 423328 555478 423337
rect 555422 423263 555478 423272
rect 555424 418192 555476 418198
rect 555424 418134 555476 418140
rect 9036 416764 9088 416770
rect 9036 416706 9088 416712
rect 9048 415449 9076 416706
rect 9034 415440 9090 415449
rect 9034 415375 9090 415384
rect 3516 404320 3568 404326
rect 3516 404262 3568 404268
rect 9404 404320 9456 404326
rect 9404 404262 9456 404268
rect 9416 403481 9444 404262
rect 9402 403472 9458 403481
rect 9402 403407 9458 403416
rect 555436 398857 555464 418134
rect 555528 411097 555556 430578
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 555514 411088 555570 411097
rect 555514 411023 555570 411032
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 555516 404388 555568 404394
rect 555516 404330 555568 404336
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 555422 398848 555478 398857
rect 555422 398783 555478 398792
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 7564 397520 7616 397526
rect 3568 397488 3570 397497
rect 7564 397462 7616 397468
rect 3514 397423 3570 397432
rect 3424 391944 3476 391950
rect 3424 391886 3476 391892
rect 3422 384432 3478 384441
rect 3422 384367 3478 384376
rect 3436 383722 3464 384367
rect 3424 383716 3476 383722
rect 3424 383658 3476 383664
rect 7576 379545 7604 397462
rect 9404 391944 9456 391950
rect 9404 391886 9456 391892
rect 9416 391513 9444 391886
rect 9402 391504 9458 391513
rect 9402 391439 9458 391448
rect 555424 390584 555476 390590
rect 555424 390526 555476 390532
rect 9036 383716 9088 383722
rect 9036 383658 9088 383664
rect 7562 379536 7618 379545
rect 7562 379471 7618 379480
rect 3422 371376 3478 371385
rect 3422 371311 3424 371320
rect 3476 371311 3478 371320
rect 8944 371340 8996 371346
rect 3424 371282 3476 371288
rect 8944 371282 8996 371288
rect 2962 358456 3018 358465
rect 2962 358391 3018 358400
rect 2976 357474 3004 358391
rect 2964 357468 3016 357474
rect 2964 357410 3016 357416
rect 6184 357468 6236 357474
rect 6184 357410 6236 357416
rect 3422 345400 3478 345409
rect 3422 345335 3424 345344
rect 3476 345335 3478 345344
rect 3424 345306 3476 345312
rect 6196 343602 6224 357410
rect 8956 355609 8984 371282
rect 9048 367577 9076 383658
rect 555436 374377 555464 390526
rect 555528 386617 555556 404330
rect 580170 391776 580226 391785
rect 580170 391711 580226 391720
rect 580184 390590 580212 391711
rect 580172 390584 580224 390590
rect 580172 390526 580224 390532
rect 555514 386608 555570 386617
rect 555514 386543 555570 386552
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 555516 378208 555568 378214
rect 555516 378150 555568 378156
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 555422 374368 555478 374377
rect 555422 374303 555478 374312
rect 9034 367568 9090 367577
rect 9034 367503 9090 367512
rect 555528 362137 555556 378150
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 555608 364404 555660 364410
rect 555608 364346 555660 364352
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 555514 362128 555570 362137
rect 555514 362063 555570 362072
rect 8942 355600 8998 355609
rect 8942 355535 8998 355544
rect 555424 351960 555476 351966
rect 555424 351902 555476 351908
rect 8944 345364 8996 345370
rect 8944 345306 8996 345312
rect 6184 343596 6236 343602
rect 6184 343538 6236 343544
rect 3422 332344 3478 332353
rect 3422 332279 3424 332288
rect 3476 332279 3478 332288
rect 7564 332308 7616 332314
rect 3424 332250 3476 332256
rect 7564 332250 7616 332256
rect 7576 319705 7604 332250
rect 8956 331673 8984 345306
rect 9402 343632 9458 343641
rect 9402 343567 9404 343576
rect 9456 343567 9458 343576
rect 9404 343538 9456 343544
rect 555436 337657 555464 351902
rect 555620 349897 555648 364346
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 555606 349888 555662 349897
rect 555606 349823 555662 349832
rect 580170 338600 580226 338609
rect 580170 338535 580226 338544
rect 580184 338162 580212 338535
rect 555516 338156 555568 338162
rect 555516 338098 555568 338104
rect 580172 338156 580224 338162
rect 580172 338098 580224 338104
rect 555422 337648 555478 337657
rect 555422 337583 555478 337592
rect 8942 331664 8998 331673
rect 8942 331599 8998 331608
rect 555528 325417 555556 338098
rect 555514 325408 555570 325417
rect 555514 325343 555570 325352
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 555424 324352 555476 324358
rect 555424 324294 555476 324300
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 7562 319696 7618 319705
rect 7562 319631 7618 319640
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 319122 3464 319223
rect 3424 319116 3476 319122
rect 3424 319058 3476 319064
rect 7656 319116 7708 319122
rect 7656 319058 7708 319064
rect 7668 307737 7696 319058
rect 555436 313177 555464 324294
rect 555422 313168 555478 313177
rect 555422 313103 555478 313112
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 555516 311908 555568 311914
rect 555516 311850 555568 311856
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 7654 307728 7710 307737
rect 7654 307663 7710 307672
rect 2778 306232 2834 306241
rect 2778 306167 2834 306176
rect 2792 305862 2820 306167
rect 2780 305856 2832 305862
rect 2780 305798 2832 305804
rect 6184 305856 6236 305862
rect 6184 305798 6236 305804
rect 6196 296682 6224 305798
rect 555528 300937 555556 311850
rect 555514 300928 555570 300937
rect 555514 300863 555570 300872
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 555424 298172 555476 298178
rect 555424 298114 555476 298120
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 6184 296676 6236 296682
rect 6184 296618 6236 296624
rect 9496 296676 9548 296682
rect 9496 296618 9548 296624
rect 9508 295769 9536 296618
rect 9494 295760 9550 295769
rect 9494 295695 9550 295704
rect 2962 293176 3018 293185
rect 2962 293111 3018 293120
rect 2976 292602 3004 293111
rect 2964 292596 3016 292602
rect 2964 292538 3016 292544
rect 6184 292596 6236 292602
rect 6184 292538 6236 292544
rect 6196 284306 6224 292538
rect 555436 288697 555464 298114
rect 555422 288688 555478 288697
rect 555422 288623 555478 288632
rect 580170 285424 580226 285433
rect 580170 285359 580226 285368
rect 580184 284374 580212 285359
rect 555424 284368 555476 284374
rect 555424 284310 555476 284316
rect 580172 284368 580224 284374
rect 580172 284310 580224 284316
rect 6184 284300 6236 284306
rect 6184 284242 6236 284248
rect 8668 284300 8720 284306
rect 8668 284242 8720 284248
rect 8680 283801 8708 284242
rect 8666 283792 8722 283801
rect 8666 283727 8722 283736
rect 3514 280120 3570 280129
rect 3514 280055 3570 280064
rect 3528 279614 3556 280055
rect 3516 279608 3568 279614
rect 3516 279550 3568 279556
rect 8208 279608 8260 279614
rect 8208 279550 8260 279556
rect 8220 271833 8248 279550
rect 555436 276457 555464 284310
rect 555422 276448 555478 276457
rect 555422 276383 555478 276392
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 555424 271924 555476 271930
rect 555424 271866 555476 271872
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 8206 271824 8262 271833
rect 8206 271759 8262 271768
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 9404 266416 9456 266422
rect 9404 266358 9456 266364
rect 9416 259865 9444 266358
rect 555436 264217 555464 271866
rect 555422 264208 555478 264217
rect 555422 264143 555478 264152
rect 9402 259856 9458 259865
rect 9402 259791 9458 259800
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 556068 258120 556120 258126
rect 556068 258062 556120 258068
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 3422 254144 3478 254153
rect 3422 254079 3424 254088
rect 3476 254079 3478 254088
rect 8944 254108 8996 254114
rect 3424 254050 3476 254056
rect 8944 254050 8996 254056
rect 8956 247897 8984 254050
rect 556080 251977 556108 258062
rect 556066 251968 556122 251977
rect 556066 251903 556122 251912
rect 8942 247888 8998 247897
rect 8942 247823 8998 247832
rect 579802 245576 579858 245585
rect 579802 245511 579858 245520
rect 579816 244322 579844 245511
rect 555424 244316 555476 244322
rect 555424 244258 555476 244264
rect 579804 244316 579856 244322
rect 579804 244258 579856 244264
rect 3698 241088 3754 241097
rect 3698 241023 3754 241032
rect 3712 235958 3740 241023
rect 555436 239737 555464 244258
rect 555422 239728 555478 239737
rect 555422 239663 555478 239672
rect 3700 235952 3752 235958
rect 9404 235952 9456 235958
rect 3700 235894 3752 235900
rect 9402 235920 9404 235929
rect 9456 235920 9458 235929
rect 9402 235855 9458 235864
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580184 231878 580212 232319
rect 555424 231872 555476 231878
rect 555424 231814 555476 231820
rect 580172 231872 580224 231878
rect 580172 231814 580224 231820
rect 4066 228032 4122 228041
rect 4122 227990 4200 228018
rect 4066 227967 4122 227976
rect 4172 224942 4200 227990
rect 555436 227497 555464 231814
rect 555422 227488 555478 227497
rect 555422 227423 555478 227432
rect 4160 224936 4212 224942
rect 4160 224878 4212 224884
rect 8852 224936 8904 224942
rect 8852 224878 8904 224884
rect 8864 223961 8892 224878
rect 8850 223952 8906 223961
rect 8850 223887 8906 223896
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 555424 218068 555476 218074
rect 555424 218010 555476 218016
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 555436 215257 555464 218010
rect 555422 215248 555478 215257
rect 555422 215183 555478 215192
rect 3146 214976 3202 214985
rect 3146 214911 3202 214920
rect 3160 213994 3188 214911
rect 3148 213988 3200 213994
rect 3148 213930 3200 213936
rect 9220 213988 9272 213994
rect 9220 213930 9272 213936
rect 9232 211993 9260 213930
rect 9218 211984 9274 211993
rect 9218 211919 9274 211928
rect 580170 205728 580226 205737
rect 555424 205692 555476 205698
rect 580170 205663 580172 205672
rect 555424 205634 555476 205640
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 555436 203017 555464 205634
rect 555422 203008 555478 203017
rect 555422 202943 555478 202952
rect 3422 201920 3478 201929
rect 3422 201855 3424 201864
rect 3476 201855 3478 201864
rect 8300 201884 8352 201890
rect 3424 201826 3476 201832
rect 8300 201826 8352 201832
rect 8312 200025 8340 201826
rect 8298 200016 8354 200025
rect 8298 199951 8354 199960
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191894 580212 192471
rect 580172 191888 580224 191894
rect 580172 191830 580224 191836
rect 555424 191820 555476 191826
rect 555424 191762 555476 191768
rect 555436 190777 555464 191762
rect 555422 190768 555478 190777
rect 555422 190703 555478 190712
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3436 188290 3464 188799
rect 3424 188284 3476 188290
rect 3424 188226 3476 188232
rect 9404 188284 9456 188290
rect 9404 188226 9456 188232
rect 9416 188057 9444 188226
rect 9402 188048 9458 188057
rect 9402 187983 9458 187992
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178702 580212 179143
rect 555424 178696 555476 178702
rect 555424 178638 555476 178644
rect 580172 178696 580224 178702
rect 580172 178638 580224 178644
rect 555436 178537 555464 178638
rect 555422 178528 555478 178537
rect 555422 178463 555478 178472
rect 9402 176080 9458 176089
rect 9402 176015 9458 176024
rect 3330 175944 3386 175953
rect 3330 175879 3386 175888
rect 3344 175642 3372 175879
rect 9416 175642 9444 176015
rect 3332 175636 3384 175642
rect 3332 175578 3384 175584
rect 9404 175636 9456 175642
rect 9404 175578 9456 175584
rect 555884 166320 555936 166326
rect 555882 166288 555884 166297
rect 580172 166320 580224 166326
rect 555936 166288 555938 166297
rect 580172 166262 580224 166268
rect 555882 166223 555938 166232
rect 580184 165889 580212 166262
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 9402 164112 9458 164121
rect 9402 164047 9458 164056
rect 9416 162926 9444 164047
rect 3424 162920 3476 162926
rect 3422 162888 3424 162897
rect 9404 162920 9456 162926
rect 3476 162888 3478 162897
rect 9404 162862 9456 162868
rect 3422 162823 3478 162832
rect 555422 154048 555478 154057
rect 555422 153983 555478 153992
rect 555436 153270 555464 153983
rect 555424 153264 555476 153270
rect 555424 153206 555476 153212
rect 579528 153264 579580 153270
rect 579528 153206 579580 153212
rect 579540 152697 579568 153206
rect 579526 152688 579582 152697
rect 579526 152623 579582 152632
rect 8206 152144 8262 152153
rect 8206 152079 8262 152088
rect 8220 150414 8248 152079
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 8208 150408 8260 150414
rect 8208 150350 8260 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 555422 141808 555478 141817
rect 555422 141743 555478 141752
rect 8206 140176 8262 140185
rect 8206 140111 8262 140120
rect 8220 137018 8248 140111
rect 555436 139398 555464 141743
rect 555424 139392 555476 139398
rect 580172 139392 580224 139398
rect 555424 139334 555476 139340
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 3240 137012 3292 137018
rect 3240 136954 3292 136960
rect 8208 137012 8260 137018
rect 8208 136954 8260 136960
rect 3252 136785 3280 136954
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 555422 129568 555478 129577
rect 555422 129503 555478 129512
rect 8206 128208 8262 128217
rect 8206 128143 8262 128152
rect 8220 123894 8248 128143
rect 555436 126954 555464 129503
rect 555424 126948 555476 126954
rect 555424 126890 555476 126896
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 3424 123888 3476 123894
rect 3424 123830 3476 123836
rect 8208 123888 8260 123894
rect 8208 123830 8260 123836
rect 3436 123729 3464 123830
rect 3422 123720 3478 123729
rect 3422 123655 3478 123664
rect 555422 117328 555478 117337
rect 555422 117263 555478 117272
rect 8942 116240 8998 116249
rect 8942 116175 8998 116184
rect 8956 110770 8984 116175
rect 555436 113150 555464 117263
rect 555424 113144 555476 113150
rect 555424 113086 555476 113092
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 3424 110764 3476 110770
rect 3424 110706 3476 110712
rect 8944 110764 8996 110770
rect 8944 110706 8996 110712
rect 3436 110673 3464 110706
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 555698 105088 555754 105097
rect 555698 105023 555754 105032
rect 9402 104272 9458 104281
rect 9402 104207 9458 104216
rect 9416 103562 9444 104207
rect 4160 103556 4212 103562
rect 4160 103498 4212 103504
rect 9404 103556 9456 103562
rect 9404 103498 9456 103504
rect 4066 97608 4122 97617
rect 4172 97594 4200 103498
rect 555712 100706 555740 105023
rect 555700 100700 555752 100706
rect 555700 100642 555752 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 4122 97566 4200 97594
rect 4066 97543 4122 97552
rect 554778 92848 554834 92857
rect 554778 92783 554834 92792
rect 9402 92304 9458 92313
rect 9402 92239 9458 92248
rect 9416 91118 9444 92239
rect 4160 91112 4212 91118
rect 4160 91054 4212 91060
rect 9404 91112 9456 91118
rect 9404 91054 9456 91060
rect 4066 84688 4122 84697
rect 4172 84674 4200 91054
rect 554792 86970 554820 92783
rect 554780 86964 554832 86970
rect 554780 86906 554832 86912
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 4122 84646 4200 84674
rect 4066 84623 4122 84632
rect 555422 80608 555478 80617
rect 555422 80543 555478 80552
rect 8942 80336 8998 80345
rect 8942 80271 8998 80280
rect 8956 71670 8984 80271
rect 555436 73166 555464 80543
rect 555424 73160 555476 73166
rect 555424 73102 555476 73108
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 3424 71664 3476 71670
rect 3422 71632 3424 71641
rect 8944 71664 8996 71670
rect 3476 71632 3478 71641
rect 8944 71606 8996 71612
rect 3422 71567 3478 71576
rect 8942 68368 8998 68377
rect 8942 68303 8998 68312
rect 555422 68368 555478 68377
rect 555422 68303 555478 68312
rect 8956 59226 8984 68303
rect 555436 60722 555464 68303
rect 555424 60716 555476 60722
rect 555424 60658 555476 60664
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 3148 59220 3200 59226
rect 3148 59162 3200 59168
rect 8944 59220 8996 59226
rect 8944 59162 8996 59168
rect 3160 58585 3188 59162
rect 3146 58576 3202 58585
rect 3146 58511 3202 58520
rect 9402 56400 9458 56409
rect 9402 56335 9458 56344
rect 9416 55282 9444 56335
rect 555422 56128 555478 56137
rect 555422 56063 555478 56072
rect 4804 55276 4856 55282
rect 4804 55218 4856 55224
rect 9404 55276 9456 55282
rect 9404 55218 9456 55224
rect 4816 45558 4844 55218
rect 555436 46918 555464 56063
rect 555424 46912 555476 46918
rect 555424 46854 555476 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 2780 45552 2832 45558
rect 2778 45520 2780 45529
rect 4804 45552 4856 45558
rect 2832 45520 2834 45529
rect 4804 45494 4856 45500
rect 2778 45455 2834 45464
rect 9402 44432 9458 44441
rect 9402 44367 9458 44376
rect 9416 44198 9444 44367
rect 3424 44192 3476 44198
rect 3424 44134 3476 44140
rect 9404 44192 9456 44198
rect 9404 44134 9456 44140
rect 3436 32473 3464 44134
rect 555422 43888 555478 43897
rect 555422 43823 555478 43832
rect 555436 33114 555464 43823
rect 580170 33144 580226 33153
rect 555424 33108 555476 33114
rect 580170 33079 580172 33088
rect 555424 33050 555476 33056
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 9402 32464 9458 32473
rect 9402 32399 9458 32408
rect 9416 31822 9444 32399
rect 3516 31816 3568 31822
rect 3516 31758 3568 31764
rect 9404 31816 9456 31822
rect 9404 31758 9456 31764
rect 3528 19417 3556 31758
rect 555514 31648 555570 31657
rect 555514 31583 555570 31592
rect 555528 20670 555556 31583
rect 555516 20664 555568 20670
rect 555516 20606 555568 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 9402 20496 9458 20505
rect 9402 20431 9458 20440
rect 3514 19408 3570 19417
rect 9416 19378 9444 20431
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 555422 19408 555478 19417
rect 3514 19343 3570 19352
rect 6184 19372 6236 19378
rect 6184 19314 6236 19320
rect 9404 19372 9456 19378
rect 555422 19343 555478 19352
rect 9404 19314 9456 19320
rect 4804 7676 4856 7682
rect 4804 7618 4856 7624
rect 3148 6520 3200 6526
rect 3146 6488 3148 6497
rect 3200 6488 3202 6497
rect 3146 6423 3202 6432
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 3052 624 3058
rect 572 2994 624 3000
rect 584 480 612 2994
rect 1688 480 1716 4830
rect 2792 3058 2820 6190
rect 4816 3534 4844 7618
rect 6196 6526 6224 19314
rect 33244 12022 33304 12050
rect 33980 12022 34316 12050
rect 34992 12022 35328 12050
rect 35912 12022 36340 12050
rect 37352 12022 37504 12050
rect 33140 9512 33192 9518
rect 33140 9454 33192 9460
rect 31300 9376 31352 9382
rect 31300 9318 31352 9324
rect 25320 9308 25372 9314
rect 25320 9250 25372 9256
rect 19432 9240 19484 9246
rect 19432 9182 19484 9188
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6184 6520 6236 6526
rect 6184 6462 6236 6468
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2884 480 2912 3470
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 480 4108 3402
rect 5264 3256 5316 3262
rect 5264 3198 5316 3204
rect 5276 480 5304 3198
rect 6472 480 6500 8910
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7668 480 7696 4762
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8772 480 8800 3606
rect 9968 480 9996 8978
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11164 480 11192 3878
rect 12360 480 12388 6122
rect 14740 3800 14792 3806
rect 14740 3742 14792 3748
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13556 480 13584 3538
rect 14752 480 14780 3742
rect 15948 480 15976 9046
rect 17040 7608 17092 7614
rect 17040 7550 17092 7556
rect 17052 480 17080 7550
rect 18236 3868 18288 3874
rect 18236 3810 18288 3816
rect 18248 480 18276 3810
rect 19444 480 19472 9182
rect 23020 9172 23072 9178
rect 23020 9114 23072 9120
rect 21824 4956 21876 4962
rect 21824 4898 21876 4904
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20640 480 20668 3674
rect 21836 480 21864 4898
rect 23032 480 23060 9114
rect 24216 4072 24268 4078
rect 24216 4014 24268 4020
rect 24228 480 24256 4014
rect 25332 480 25360 9250
rect 30104 7744 30156 7750
rect 30104 7686 30156 7692
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 26528 480 26556 6258
rect 28908 4004 28960 4010
rect 28908 3946 28960 3952
rect 27712 3324 27764 3330
rect 27712 3266 27764 3272
rect 27724 480 27752 3266
rect 28920 480 28948 3946
rect 30116 480 30144 7686
rect 31312 480 31340 9318
rect 33152 4894 33180 9454
rect 33244 6254 33272 12022
rect 33980 9518 34008 12022
rect 33968 9512 34020 9518
rect 33968 9454 34020 9460
rect 34992 7682 35020 12022
rect 34980 7676 35032 7682
rect 34980 7618 35032 7624
rect 33232 6248 33284 6254
rect 33232 6190 33284 6196
rect 33140 4888 33192 4894
rect 33140 4830 33192 4836
rect 33600 4888 33652 4894
rect 33600 4830 33652 4836
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 32416 480 32444 3062
rect 33612 480 33640 4830
rect 34796 4140 34848 4146
rect 34796 4082 34848 4088
rect 34808 480 34836 4082
rect 35912 3534 35940 12022
rect 37188 6248 37240 6254
rect 37188 6190 37240 6196
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 36004 480 36032 3470
rect 37200 480 37228 6190
rect 37476 3262 37504 12022
rect 38028 12022 38364 12050
rect 38672 12022 39376 12050
rect 40236 12022 40388 12050
rect 41064 12022 41400 12050
rect 41708 12022 42412 12050
rect 42812 12022 43424 12050
rect 44376 12022 44436 12050
rect 45112 12022 45448 12050
rect 46124 12022 46460 12050
rect 47136 12022 47472 12050
rect 38028 8974 38056 12022
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 38672 4826 38700 12022
rect 38660 4820 38712 4826
rect 38660 4762 38712 4768
rect 40236 3670 40264 12022
rect 41064 9042 41092 12022
rect 41052 9036 41104 9042
rect 41052 8978 41104 8984
rect 41708 6914 41736 12022
rect 41432 6886 41736 6914
rect 40684 4820 40736 4826
rect 40684 4762 40736 4768
rect 40224 3664 40276 3670
rect 40224 3606 40276 3612
rect 38384 3460 38436 3466
rect 38384 3402 38436 3408
rect 37464 3256 37516 3262
rect 37464 3198 37516 3204
rect 38396 480 38424 3402
rect 39578 3360 39634 3369
rect 39578 3295 39634 3304
rect 39592 480 39620 3295
rect 40696 480 40724 4762
rect 41432 3942 41460 6886
rect 42812 6186 42840 12022
rect 44180 9512 44232 9518
rect 44180 9454 44232 9460
rect 42800 6180 42852 6186
rect 42800 6122 42852 6128
rect 41420 3936 41472 3942
rect 41420 3878 41472 3884
rect 41880 3936 41932 3942
rect 41880 3878 41932 3884
rect 41892 480 41920 3878
rect 44192 3806 44220 9454
rect 44180 3800 44232 3806
rect 44180 3742 44232 3748
rect 44272 3800 44324 3806
rect 44272 3742 44324 3748
rect 43076 3664 43128 3670
rect 43076 3606 43128 3612
rect 43088 480 43116 3606
rect 44284 480 44312 3742
rect 44376 3602 44404 12022
rect 45112 9518 45140 12022
rect 45100 9512 45152 9518
rect 45100 9454 45152 9460
rect 46124 9110 46152 12022
rect 46112 9104 46164 9110
rect 46112 9046 46164 9052
rect 47136 7614 47164 12022
rect 48470 11778 48498 12036
rect 49160 12022 49496 12050
rect 49804 12022 50508 12050
rect 51092 12022 51520 12050
rect 52472 12022 52532 12050
rect 52656 12022 53544 12050
rect 54220 12022 54556 12050
rect 55324 12022 55568 12050
rect 56244 12022 56580 12050
rect 56704 12022 57592 12050
rect 58268 12022 58604 12050
rect 59372 12022 59616 12050
rect 59832 12022 60628 12050
rect 60752 12022 61640 12050
rect 62132 12022 62652 12050
rect 63604 12022 63664 12050
rect 64340 12022 64676 12050
rect 64892 12022 65688 12050
rect 66272 12022 66700 12050
rect 48470 11750 48544 11778
rect 47860 7812 47912 7818
rect 47860 7754 47912 7760
rect 47124 7608 47176 7614
rect 47124 7550 47176 7556
rect 44364 3596 44416 3602
rect 44364 3538 44416 3544
rect 46664 3596 46716 3602
rect 46664 3538 46716 3544
rect 45468 3256 45520 3262
rect 45468 3198 45520 3204
rect 45480 480 45508 3198
rect 46676 480 46704 3538
rect 47872 480 47900 7754
rect 48516 3874 48544 11750
rect 49160 9246 49188 12022
rect 49148 9240 49200 9246
rect 49148 9182 49200 9188
rect 48504 3868 48556 3874
rect 48504 3810 48556 3816
rect 49804 3738 49832 12022
rect 50160 8968 50212 8974
rect 50160 8910 50212 8916
rect 49792 3732 49844 3738
rect 49792 3674 49844 3680
rect 48964 3052 49016 3058
rect 48964 2994 49016 3000
rect 48976 480 49004 2994
rect 50172 480 50200 8910
rect 51092 4962 51120 12022
rect 52472 9178 52500 12022
rect 52460 9172 52512 9178
rect 52460 9114 52512 9120
rect 52656 6914 52684 12022
rect 54220 9314 54248 12022
rect 55220 9512 55272 9518
rect 55220 9454 55272 9460
rect 54208 9308 54260 9314
rect 54208 9250 54260 9256
rect 52564 6886 52684 6914
rect 51080 4956 51132 4962
rect 51080 4898 51132 4904
rect 51356 4956 51408 4962
rect 51356 4898 51408 4904
rect 51368 480 51396 4898
rect 52564 4078 52592 6886
rect 54944 6180 54996 6186
rect 54944 6122 54996 6128
rect 52552 4072 52604 4078
rect 52552 4014 52604 4020
rect 53748 3732 53800 3738
rect 53748 3674 53800 3680
rect 52552 3188 52604 3194
rect 52552 3130 52604 3136
rect 52564 480 52592 3130
rect 53760 480 53788 3674
rect 54956 480 54984 6122
rect 55232 3330 55260 9454
rect 55324 6322 55352 12022
rect 56244 9518 56272 12022
rect 56232 9512 56284 9518
rect 56232 9454 56284 9460
rect 55312 6316 55364 6322
rect 55312 6258 55364 6264
rect 56048 4072 56100 4078
rect 56048 4014 56100 4020
rect 55220 3324 55272 3330
rect 55220 3266 55272 3272
rect 56060 480 56088 4014
rect 56704 4010 56732 12022
rect 57244 9036 57296 9042
rect 57244 8978 57296 8984
rect 56692 4004 56744 4010
rect 56692 3946 56744 3952
rect 57256 480 57284 8978
rect 58268 7750 58296 12022
rect 59372 9382 59400 12022
rect 59360 9376 59412 9382
rect 59360 9318 59412 9324
rect 58256 7744 58308 7750
rect 58256 7686 58308 7692
rect 58440 7608 58492 7614
rect 58440 7550 58492 7556
rect 58452 480 58480 7550
rect 59832 6914 59860 12022
rect 59556 6886 59860 6914
rect 59556 3126 59584 6886
rect 60752 4894 60780 12022
rect 60740 4888 60792 4894
rect 60740 4830 60792 4836
rect 62028 4888 62080 4894
rect 62028 4830 62080 4836
rect 60832 4004 60884 4010
rect 60832 3946 60884 3952
rect 59636 3392 59688 3398
rect 59636 3334 59688 3340
rect 59544 3120 59596 3126
rect 59544 3062 59596 3068
rect 59648 480 59676 3334
rect 60844 480 60872 3946
rect 62040 480 62068 4830
rect 62132 4146 62160 12022
rect 63408 9444 63460 9450
rect 63408 9386 63460 9392
rect 63420 6254 63448 9386
rect 63408 6248 63460 6254
rect 63408 6190 63460 6196
rect 62120 4140 62172 4146
rect 62120 4082 62172 4088
rect 63224 4140 63276 4146
rect 63224 4082 63276 4088
rect 63236 480 63264 4082
rect 63604 3534 63632 12022
rect 64340 9450 64368 12022
rect 64328 9444 64380 9450
rect 64328 9386 64380 9392
rect 64328 9104 64380 9110
rect 64328 9046 64380 9052
rect 63592 3528 63644 3534
rect 63592 3470 63644 3476
rect 64340 480 64368 9046
rect 64892 3466 64920 12022
rect 65524 6248 65576 6254
rect 65524 6190 65576 6196
rect 64880 3460 64932 3466
rect 64880 3402 64932 3408
rect 65536 480 65564 6190
rect 66272 3369 66300 12022
rect 67698 11778 67726 12036
rect 68388 12022 68724 12050
rect 69032 12022 69736 12050
rect 70504 12022 70748 12050
rect 71424 12022 71760 12050
rect 71884 12022 72772 12050
rect 73448 12022 73784 12050
rect 74736 12022 74796 12050
rect 75472 12022 75808 12050
rect 75932 12022 76820 12050
rect 77312 12022 77832 12050
rect 78692 12022 78844 12050
rect 78968 12022 79856 12050
rect 80072 12022 80868 12050
rect 81544 12022 81880 12050
rect 82832 12022 82892 12050
rect 83108 12022 83904 12050
rect 84212 12022 84916 12050
rect 85684 12022 85928 12050
rect 86604 12022 86940 12050
rect 87616 12022 87952 12050
rect 88352 12022 88964 12050
rect 89824 12022 89976 12050
rect 90652 12022 90988 12050
rect 91664 12022 92000 12050
rect 92584 12022 93012 12050
rect 93964 12022 94024 12050
rect 94700 12022 95036 12050
rect 95252 12022 96048 12050
rect 96632 12022 97060 12050
rect 67698 11750 67772 11778
rect 67640 9512 67692 9518
rect 67640 9454 67692 9460
rect 67652 3942 67680 9454
rect 67744 4826 67772 11750
rect 68388 9518 68416 12022
rect 68376 9512 68428 9518
rect 68376 9454 68428 9460
rect 67732 4820 67784 4826
rect 67732 4762 67784 4768
rect 67640 3936 67692 3942
rect 67640 3878 67692 3884
rect 67916 3936 67968 3942
rect 67916 3878 67968 3884
rect 66720 3460 66772 3466
rect 66720 3402 66772 3408
rect 66258 3360 66314 3369
rect 66258 3295 66314 3304
rect 66732 480 66760 3402
rect 67928 480 67956 3878
rect 69032 3670 69060 12022
rect 70400 9512 70452 9518
rect 70400 9454 70452 9460
rect 69112 7676 69164 7682
rect 69112 7618 69164 7624
rect 69020 3664 69072 3670
rect 69020 3606 69072 3612
rect 69124 480 69152 7618
rect 70308 3528 70360 3534
rect 70308 3470 70360 3476
rect 70320 480 70348 3470
rect 70412 3262 70440 9454
rect 70504 3806 70532 12022
rect 71424 9518 71452 12022
rect 71412 9512 71464 9518
rect 71412 9454 71464 9460
rect 71884 6914 71912 12022
rect 73448 7818 73476 12022
rect 73436 7812 73488 7818
rect 73436 7754 73488 7760
rect 71792 6886 71912 6914
rect 70492 3800 70544 3806
rect 70492 3742 70544 3748
rect 71504 3664 71556 3670
rect 71504 3606 71556 3612
rect 70400 3256 70452 3262
rect 70400 3198 70452 3204
rect 71516 480 71544 3606
rect 71792 3602 71820 6886
rect 72608 5024 72660 5030
rect 72608 4966 72660 4972
rect 71780 3596 71832 3602
rect 71780 3538 71832 3544
rect 72620 480 72648 4966
rect 73804 3596 73856 3602
rect 73804 3538 73856 3544
rect 73816 480 73844 3538
rect 74736 3058 74764 12022
rect 75472 8974 75500 12022
rect 75460 8968 75512 8974
rect 75460 8910 75512 8916
rect 75932 4962 75960 12022
rect 76196 6316 76248 6322
rect 76196 6258 76248 6264
rect 75920 4956 75972 4962
rect 75920 4898 75972 4904
rect 75000 3800 75052 3806
rect 75000 3742 75052 3748
rect 74724 3052 74776 3058
rect 74724 2994 74776 3000
rect 75012 480 75040 3742
rect 76208 480 76236 6258
rect 77312 3194 77340 12022
rect 78692 3738 78720 12022
rect 78968 6914 78996 12022
rect 78784 6886 78996 6914
rect 78784 6186 78812 6886
rect 78772 6180 78824 6186
rect 78772 6122 78824 6128
rect 79692 4820 79744 4826
rect 79692 4762 79744 4768
rect 78680 3732 78732 3738
rect 78680 3674 78732 3680
rect 78586 3360 78642 3369
rect 77392 3324 77444 3330
rect 78586 3295 78642 3304
rect 77392 3266 77444 3272
rect 77300 3188 77352 3194
rect 77300 3130 77352 3136
rect 77404 480 77432 3266
rect 78600 480 78628 3295
rect 79704 480 79732 4762
rect 80072 4078 80100 12022
rect 81544 9042 81572 12022
rect 81532 9036 81584 9042
rect 81532 8978 81584 8984
rect 82832 7614 82860 12022
rect 82820 7608 82872 7614
rect 82820 7550 82872 7556
rect 83108 6914 83136 12022
rect 82832 6886 83136 6914
rect 80060 4072 80112 4078
rect 80060 4014 80112 4020
rect 82832 3398 82860 6886
rect 84212 4010 84240 12022
rect 85580 9512 85632 9518
rect 85580 9454 85632 9460
rect 85592 4146 85620 9454
rect 85684 4894 85712 12022
rect 86604 9518 86632 12022
rect 86592 9512 86644 9518
rect 86592 9454 86644 9460
rect 87616 9110 87644 12022
rect 87604 9104 87656 9110
rect 87604 9046 87656 9052
rect 87420 8356 87472 8362
rect 87420 8298 87472 8304
rect 87432 5030 87460 8298
rect 88352 6254 88380 12022
rect 89720 9512 89772 9518
rect 89720 9454 89772 9460
rect 88524 9240 88576 9246
rect 88524 9182 88576 9188
rect 88340 6248 88392 6254
rect 88340 6190 88392 6196
rect 87420 5024 87472 5030
rect 87420 4966 87472 4972
rect 85672 4888 85724 4894
rect 85672 4830 85724 4836
rect 85580 4140 85632 4146
rect 85580 4082 85632 4088
rect 85672 4072 85724 4078
rect 85672 4014 85724 4020
rect 84200 4004 84252 4010
rect 84200 3946 84252 3952
rect 84476 3732 84528 3738
rect 84476 3674 84528 3680
rect 82820 3392 82872 3398
rect 82820 3334 82872 3340
rect 83280 3392 83332 3398
rect 83280 3334 83332 3340
rect 80888 3256 80940 3262
rect 80888 3198 80940 3204
rect 80900 480 80928 3198
rect 82084 3188 82136 3194
rect 82084 3130 82136 3136
rect 82096 480 82124 3130
rect 83292 480 83320 3334
rect 84488 480 84516 3674
rect 85684 480 85712 4014
rect 86868 4004 86920 4010
rect 86868 3946 86920 3952
rect 86880 480 86908 3946
rect 87972 3868 88024 3874
rect 87972 3810 88024 3816
rect 87984 480 88012 3810
rect 88536 3194 88564 9182
rect 88892 9172 88944 9178
rect 88892 9114 88944 9120
rect 88904 3398 88932 9114
rect 89168 4140 89220 4146
rect 89168 4082 89220 4088
rect 88892 3392 88944 3398
rect 88892 3334 88944 3340
rect 88524 3188 88576 3194
rect 88524 3130 88576 3136
rect 89180 480 89208 4082
rect 89732 3942 89760 9454
rect 89720 3936 89772 3942
rect 89720 3878 89772 3884
rect 89824 3466 89852 12022
rect 90652 9518 90680 12022
rect 90640 9512 90692 9518
rect 90640 9454 90692 9460
rect 91664 7682 91692 12022
rect 91652 7676 91704 7682
rect 91652 7618 91704 7624
rect 90364 3936 90416 3942
rect 90364 3878 90416 3884
rect 89812 3460 89864 3466
rect 89812 3402 89864 3408
rect 90376 480 90404 3878
rect 92584 3534 92612 12022
rect 92756 8968 92808 8974
rect 92756 8910 92808 8916
rect 92572 3528 92624 3534
rect 92572 3470 92624 3476
rect 91560 3460 91612 3466
rect 91560 3402 91612 3408
rect 91572 480 91600 3402
rect 92768 480 92796 8910
rect 93964 3670 93992 12022
rect 94700 8362 94728 12022
rect 94688 8356 94740 8362
rect 94688 8298 94740 8304
rect 93952 3664 94004 3670
rect 93952 3606 94004 3612
rect 95252 3602 95280 12022
rect 96632 3806 96660 12022
rect 98058 11778 98086 12036
rect 98748 12022 99084 12050
rect 99760 12022 100096 12050
rect 100772 12022 101108 12050
rect 101784 12022 102120 12050
rect 102796 12022 103132 12050
rect 103808 12022 104144 12050
rect 104912 12022 105156 12050
rect 105832 12022 106168 12050
rect 106844 12022 107180 12050
rect 107856 12022 108192 12050
rect 109052 12022 109204 12050
rect 109880 12022 110216 12050
rect 110892 12022 111228 12050
rect 111812 12022 112240 12050
rect 113192 12022 113252 12050
rect 113928 12022 114264 12050
rect 114940 12022 115276 12050
rect 115952 12022 116288 12050
rect 117056 12022 117300 12050
rect 117976 12022 118312 12050
rect 118712 12022 119324 12050
rect 120092 12022 120336 12050
rect 121012 12022 121348 12050
rect 122024 12022 122360 12050
rect 123036 12022 123372 12050
rect 124232 12022 124384 12050
rect 124784 12022 125396 12050
rect 125612 12022 126408 12050
rect 126992 12022 127420 12050
rect 128372 12022 128432 12050
rect 129108 12022 129444 12050
rect 129752 12022 130456 12050
rect 131316 12022 131468 12050
rect 132144 12022 132480 12050
rect 132604 12022 133492 12050
rect 134168 12022 134504 12050
rect 98058 11750 98132 11778
rect 97908 9444 97960 9450
rect 97908 9386 97960 9392
rect 96620 3800 96672 3806
rect 96620 3742 96672 3748
rect 97448 3800 97500 3806
rect 97448 3742 97500 3748
rect 96252 3664 96304 3670
rect 96252 3606 96304 3612
rect 95240 3596 95292 3602
rect 95240 3538 95292 3544
rect 93952 3392 94004 3398
rect 93952 3334 94004 3340
rect 93964 480 93992 3334
rect 95148 3188 95200 3194
rect 95148 3130 95200 3136
rect 95160 480 95188 3130
rect 96264 480 96292 3606
rect 97460 480 97488 3742
rect 97920 3330 97948 9386
rect 98104 6322 98132 11750
rect 98748 9450 98776 12022
rect 98736 9444 98788 9450
rect 98736 9386 98788 9392
rect 98552 9104 98604 9110
rect 98552 9046 98604 9052
rect 98092 6316 98144 6322
rect 98092 6258 98144 6264
rect 97908 3324 97960 3330
rect 97908 3266 97960 3272
rect 98564 3262 98592 9046
rect 99760 3369 99788 12022
rect 99840 9036 99892 9042
rect 99840 8978 99892 8984
rect 99746 3360 99802 3369
rect 99746 3295 99802 3304
rect 98552 3256 98604 3262
rect 98552 3198 98604 3204
rect 98644 3120 98696 3126
rect 98644 3062 98696 3068
rect 98656 480 98684 3062
rect 99852 480 99880 8978
rect 100772 4826 100800 12022
rect 101784 9110 101812 12022
rect 102796 9246 102824 12022
rect 102784 9240 102836 9246
rect 102784 9182 102836 9188
rect 103808 9178 103836 12022
rect 103796 9172 103848 9178
rect 103796 9114 103848 9120
rect 103980 9172 104032 9178
rect 103980 9114 104032 9120
rect 101772 9104 101824 9110
rect 101772 9046 101824 9052
rect 103336 9104 103388 9110
rect 103336 9046 103388 9052
rect 100760 4820 100812 4826
rect 100760 4762 100812 4768
rect 101876 3998 102088 4026
rect 101876 3738 101904 3998
rect 102060 3874 102088 3998
rect 101956 3868 102008 3874
rect 101956 3810 102008 3816
rect 102048 3868 102100 3874
rect 102048 3810 102100 3816
rect 101864 3732 101916 3738
rect 101864 3674 101916 3680
rect 101036 3528 101088 3534
rect 101036 3470 101088 3476
rect 101048 480 101076 3470
rect 101968 3262 101996 3810
rect 102232 3324 102284 3330
rect 102232 3266 102284 3272
rect 101956 3256 102008 3262
rect 101956 3198 102008 3204
rect 102244 480 102272 3266
rect 103348 480 103376 9046
rect 103992 3670 104020 9114
rect 104912 3874 104940 12022
rect 105832 4078 105860 12022
rect 106280 8832 106332 8838
rect 106280 8774 106332 8780
rect 106292 4146 106320 8774
rect 106280 4140 106332 4146
rect 106280 4082 106332 4088
rect 105820 4072 105872 4078
rect 105820 4014 105872 4020
rect 106844 4010 106872 12022
rect 107660 9512 107712 9518
rect 107660 9454 107712 9460
rect 106832 4004 106884 4010
rect 106832 3946 106884 3952
rect 107672 3942 107700 9454
rect 107660 3936 107712 3942
rect 107660 3878 107712 3884
rect 104900 3868 104952 3874
rect 104900 3810 104952 3816
rect 103980 3664 104032 3670
rect 103980 3606 104032 3612
rect 106924 3664 106976 3670
rect 106924 3606 106976 3612
rect 104624 3596 104676 3602
rect 104624 3538 104676 3544
rect 104636 1850 104664 3538
rect 105728 3392 105780 3398
rect 105728 3334 105780 3340
rect 104544 1822 104664 1850
rect 104544 480 104572 1822
rect 105740 480 105768 3334
rect 106936 480 106964 3606
rect 107856 3262 107884 12022
rect 109052 8838 109080 12022
rect 109880 9518 109908 12022
rect 110892 9518 110920 12022
rect 109868 9512 109920 9518
rect 109868 9454 109920 9460
rect 110328 9512 110380 9518
rect 110328 9454 110380 9460
rect 110880 9512 110932 9518
rect 110880 9454 110932 9460
rect 109040 8832 109092 8838
rect 109040 8774 109092 8780
rect 109776 8424 109828 8430
rect 109776 8366 109828 8372
rect 109684 8356 109736 8362
rect 109684 8298 109736 8304
rect 108120 4004 108172 4010
rect 108120 3946 108172 3952
rect 107844 3256 107896 3262
rect 107844 3198 107896 3204
rect 108132 480 108160 3946
rect 109316 3868 109368 3874
rect 109316 3810 109368 3816
rect 109328 480 109356 3810
rect 109696 3466 109724 8298
rect 109684 3460 109736 3466
rect 109684 3402 109736 3408
rect 109788 3194 109816 8366
rect 110340 3738 110368 9454
rect 111064 9240 111116 9246
rect 111064 9182 111116 9188
rect 110512 3936 110564 3942
rect 110512 3878 110564 3884
rect 110328 3732 110380 3738
rect 110328 3674 110380 3680
rect 109776 3188 109828 3194
rect 109776 3130 109828 3136
rect 110524 480 110552 3878
rect 111076 3126 111104 9182
rect 111812 8974 111840 12022
rect 111984 9376 112036 9382
rect 111984 9318 112036 9324
rect 111800 8968 111852 8974
rect 111800 8910 111852 8916
rect 111892 8968 111944 8974
rect 111892 8910 111944 8916
rect 111616 3460 111668 3466
rect 111616 3402 111668 3408
rect 111064 3120 111116 3126
rect 111064 3062 111116 3068
rect 111628 480 111656 3402
rect 111904 3398 111932 8910
rect 111996 3806 112024 9318
rect 113192 8362 113220 12022
rect 113928 8430 113956 12022
rect 114940 9178 114968 12022
rect 115952 9382 115980 12022
rect 116952 9512 117004 9518
rect 116952 9454 117004 9460
rect 115940 9376 115992 9382
rect 115940 9318 115992 9324
rect 114928 9172 114980 9178
rect 114928 9114 114980 9120
rect 113916 8424 113968 8430
rect 113916 8366 113968 8372
rect 113180 8356 113232 8362
rect 113180 8298 113232 8304
rect 116400 4140 116452 4146
rect 116400 4082 116452 4088
rect 111984 3800 112036 3806
rect 111984 3742 112036 3748
rect 115204 3800 115256 3806
rect 115204 3742 115256 3748
rect 114008 3732 114060 3738
rect 114008 3674 114060 3680
rect 111892 3392 111944 3398
rect 111892 3334 111944 3340
rect 112812 3392 112864 3398
rect 112812 3334 112864 3340
rect 112824 480 112852 3334
rect 114020 480 114048 3674
rect 115216 480 115244 3742
rect 116412 480 116440 4082
rect 116964 3330 116992 9454
rect 117056 9246 117084 12022
rect 117044 9240 117096 9246
rect 117044 9182 117096 9188
rect 117976 9042 118004 12022
rect 117964 9036 118016 9042
rect 117964 8978 118016 8984
rect 117596 4072 117648 4078
rect 117596 4014 117648 4020
rect 116952 3324 117004 3330
rect 116952 3266 117004 3272
rect 117608 480 117636 4014
rect 118712 3534 118740 12022
rect 120092 9518 120120 12022
rect 120080 9512 120132 9518
rect 120080 9454 120132 9460
rect 121012 9110 121040 12022
rect 122024 9518 122052 12022
rect 121368 9512 121420 9518
rect 121368 9454 121420 9460
rect 122012 9512 122064 9518
rect 122012 9454 122064 9460
rect 121000 9104 121052 9110
rect 121000 9046 121052 9052
rect 121380 3602 121408 9454
rect 123036 8974 123064 12022
rect 124232 9466 124260 12022
rect 124140 9438 124260 9466
rect 123024 8968 123076 8974
rect 123024 8910 123076 8916
rect 124140 3670 124168 9438
rect 124784 6914 124812 12022
rect 124324 6886 124812 6914
rect 124324 4010 124352 6886
rect 124312 4004 124364 4010
rect 124312 3946 124364 3952
rect 125612 3874 125640 12022
rect 126888 9376 126940 9382
rect 126888 9318 126940 9324
rect 126244 8628 126296 8634
rect 126244 8570 126296 8576
rect 125600 3868 125652 3874
rect 125600 3810 125652 3816
rect 125876 3868 125928 3874
rect 125876 3810 125928 3816
rect 124128 3664 124180 3670
rect 124128 3606 124180 3612
rect 121368 3596 121420 3602
rect 121368 3538 121420 3544
rect 118700 3528 118752 3534
rect 118700 3470 118752 3476
rect 119896 3528 119948 3534
rect 119896 3470 119948 3476
rect 118792 3188 118844 3194
rect 118792 3130 118844 3136
rect 118804 480 118832 3130
rect 119908 480 119936 3470
rect 121092 3324 121144 3330
rect 121092 3266 121144 3272
rect 121104 480 121132 3266
rect 122288 3256 122340 3262
rect 122288 3198 122340 3204
rect 124680 3256 124732 3262
rect 124680 3198 124732 3204
rect 122300 480 122328 3198
rect 123484 3052 123536 3058
rect 123484 2994 123536 3000
rect 123496 480 123524 2994
rect 124692 480 124720 3198
rect 125888 480 125916 3810
rect 126256 3398 126284 8570
rect 126244 3392 126296 3398
rect 126244 3334 126296 3340
rect 126900 2990 126928 9318
rect 126992 3942 127020 12022
rect 128372 9466 128400 12022
rect 128280 9438 128400 9466
rect 127164 9172 127216 9178
rect 127164 9114 127216 9120
rect 126980 3936 127032 3942
rect 126980 3878 127032 3884
rect 126980 3392 127032 3398
rect 126980 3334 127032 3340
rect 126888 2984 126940 2990
rect 126888 2926 126940 2932
rect 126992 480 127020 3334
rect 127176 3330 127204 9114
rect 128176 4004 128228 4010
rect 128176 3946 128228 3952
rect 127164 3324 127216 3330
rect 127164 3266 127216 3272
rect 128188 480 128216 3946
rect 128280 3466 128308 9438
rect 129108 8634 129136 12022
rect 129648 8968 129700 8974
rect 129648 8910 129700 8916
rect 129096 8628 129148 8634
rect 129096 8570 129148 8576
rect 128268 3460 128320 3466
rect 128268 3402 128320 3408
rect 129372 3460 129424 3466
rect 129372 3402 129424 3408
rect 129384 480 129412 3402
rect 129660 3126 129688 8910
rect 129752 3738 129780 12022
rect 131028 9512 131080 9518
rect 131028 9454 131080 9460
rect 130384 9240 130436 9246
rect 130384 9182 130436 9188
rect 129740 3732 129792 3738
rect 129740 3674 129792 3680
rect 129648 3120 129700 3126
rect 129648 3062 129700 3068
rect 130396 3058 130424 9182
rect 131040 4146 131068 9454
rect 131120 9104 131172 9110
rect 131120 9046 131172 9052
rect 131028 4140 131080 4146
rect 131028 4082 131080 4088
rect 130568 3732 130620 3738
rect 130568 3674 130620 3680
rect 130384 3052 130436 3058
rect 130384 2994 130436 3000
rect 130580 480 130608 3674
rect 131132 3262 131160 9046
rect 131316 3806 131344 12022
rect 132144 9518 132172 12022
rect 132132 9512 132184 9518
rect 132604 9466 132632 12022
rect 132132 9454 132184 9460
rect 132512 9438 132632 9466
rect 133972 9512 134024 9518
rect 133972 9454 134024 9460
rect 131764 4140 131816 4146
rect 131764 4082 131816 4088
rect 131304 3800 131356 3806
rect 131304 3742 131356 3748
rect 131120 3256 131172 3262
rect 131120 3198 131172 3204
rect 131776 480 131804 4082
rect 132512 4078 132540 9438
rect 132592 9308 132644 9314
rect 132592 9250 132644 9256
rect 132500 4072 132552 4078
rect 132500 4014 132552 4020
rect 132604 3874 132632 9250
rect 133880 9036 133932 9042
rect 133880 8978 133932 8984
rect 133892 4010 133920 8978
rect 133880 4004 133932 4010
rect 133880 3946 133932 3952
rect 132592 3868 132644 3874
rect 132592 3810 132644 3816
rect 132960 3868 133012 3874
rect 132960 3810 133012 3816
rect 132972 480 133000 3810
rect 133984 3398 134012 9454
rect 134168 9382 134196 12022
rect 135502 11778 135530 12036
rect 136192 12022 136528 12050
rect 137204 12022 137540 12050
rect 138216 12022 138552 12050
rect 139412 12022 139564 12050
rect 140240 12022 140576 12050
rect 141252 12022 141588 12050
rect 142356 12022 142600 12050
rect 143552 12022 143612 12050
rect 144288 12022 144624 12050
rect 145300 12022 145636 12050
rect 146312 12022 146648 12050
rect 147324 12022 147660 12050
rect 148336 12022 148672 12050
rect 149348 12022 149684 12050
rect 150452 12022 150696 12050
rect 151372 12022 151708 12050
rect 152384 12022 152720 12050
rect 153396 12022 153732 12050
rect 154592 12022 154744 12050
rect 155420 12022 155756 12050
rect 156432 12022 156768 12050
rect 157444 12022 157780 12050
rect 158732 12022 158792 12050
rect 159468 12022 159804 12050
rect 160480 12022 160816 12050
rect 161676 12022 161828 12050
rect 162504 12022 162840 12050
rect 163516 12022 163852 12050
rect 164528 12022 164864 12050
rect 165632 12022 165876 12050
rect 166552 12022 166888 12050
rect 167564 12022 167900 12050
rect 168576 12022 168912 12050
rect 169772 12022 169924 12050
rect 170600 12022 170936 12050
rect 171612 12022 171948 12050
rect 172624 12022 172960 12050
rect 173912 12022 173972 12050
rect 174648 12022 174984 12050
rect 175660 12022 175996 12050
rect 176672 12022 177008 12050
rect 177684 12022 178020 12050
rect 178696 12022 179032 12050
rect 179432 12022 180044 12050
rect 180812 12022 181056 12050
rect 181272 12022 182068 12050
rect 182192 12022 183080 12050
rect 183572 12022 184092 12050
rect 184952 12022 185104 12050
rect 185228 12022 186116 12050
rect 186332 12022 187128 12050
rect 187712 12022 188140 12050
rect 189092 12022 189152 12050
rect 189368 12022 190164 12050
rect 190472 12022 191176 12050
rect 191852 12022 192188 12050
rect 192312 12022 193200 12050
rect 193508 12022 194212 12050
rect 194612 12022 195224 12050
rect 195992 12022 196236 12050
rect 196360 12022 197248 12050
rect 197372 12022 198260 12050
rect 198752 12022 199272 12050
rect 200224 12022 200284 12050
rect 200960 12022 201296 12050
rect 201604 12022 202308 12050
rect 202892 12022 203320 12050
rect 135502 11750 135576 11778
rect 134156 9376 134208 9382
rect 134156 9318 134208 9324
rect 135260 3936 135312 3942
rect 135260 3878 135312 3884
rect 133972 3392 134024 3398
rect 133972 3334 134024 3340
rect 134156 2984 134208 2990
rect 134156 2926 134208 2932
rect 134168 480 134196 2926
rect 135272 480 135300 3878
rect 135548 3534 135576 11750
rect 136192 9178 136220 12022
rect 136180 9172 136232 9178
rect 136180 9114 136232 9120
rect 136548 9172 136600 9178
rect 136548 9114 136600 9120
rect 136456 4072 136508 4078
rect 136456 4014 136508 4020
rect 135536 3528 135588 3534
rect 135536 3470 135588 3476
rect 136468 480 136496 4014
rect 136560 3466 136588 9114
rect 137204 8974 137232 12022
rect 138216 9246 138244 12022
rect 138204 9240 138256 9246
rect 138204 9182 138256 9188
rect 139412 9110 139440 12022
rect 140240 9314 140268 12022
rect 141252 9518 141280 12022
rect 141240 9512 141292 9518
rect 141240 9454 141292 9460
rect 140872 9444 140924 9450
rect 140872 9386 140924 9392
rect 140228 9308 140280 9314
rect 140228 9250 140280 9256
rect 140044 9240 140096 9246
rect 140044 9182 140096 9188
rect 139400 9104 139452 9110
rect 139400 9046 139452 9052
rect 137192 8968 137244 8974
rect 137192 8910 137244 8916
rect 138204 8968 138256 8974
rect 138204 8910 138256 8916
rect 137100 8356 137152 8362
rect 137100 8298 137152 8304
rect 137112 3738 137140 8298
rect 138216 4146 138244 8910
rect 138204 4140 138256 4146
rect 138204 4082 138256 4088
rect 137652 4004 137704 4010
rect 137652 3946 137704 3952
rect 137100 3732 137152 3738
rect 137100 3674 137152 3680
rect 136548 3460 136600 3466
rect 136548 3402 136600 3408
rect 137664 480 137692 3946
rect 140056 3874 140084 9182
rect 140044 3868 140096 3874
rect 140044 3810 140096 3816
rect 138848 3800 138900 3806
rect 138848 3742 138900 3748
rect 138860 480 138888 3742
rect 140044 3732 140096 3738
rect 140044 3674 140096 3680
rect 140056 480 140084 3674
rect 140884 2990 140912 9386
rect 142252 9376 142304 9382
rect 142252 9318 142304 9324
rect 142264 4078 142292 9318
rect 142356 9042 142384 12022
rect 143552 9178 143580 12022
rect 143632 9580 143684 9586
rect 143632 9522 143684 9528
rect 143540 9172 143592 9178
rect 143540 9114 143592 9120
rect 142344 9036 142396 9042
rect 142344 8978 142396 8984
rect 142344 8900 142396 8906
rect 142344 8842 142396 8848
rect 142252 4072 142304 4078
rect 142252 4014 142304 4020
rect 142356 3942 142384 8842
rect 143644 4010 143672 9522
rect 144288 8362 144316 12022
rect 145300 8974 145328 12022
rect 146208 9512 146260 9518
rect 146208 9454 146260 9460
rect 145288 8968 145340 8974
rect 145288 8910 145340 8916
rect 144276 8356 144328 8362
rect 144276 8298 144328 8304
rect 143632 4004 143684 4010
rect 143632 3946 143684 3952
rect 142344 3936 142396 3942
rect 142344 3878 142396 3884
rect 141240 3868 141292 3874
rect 141240 3810 141292 3816
rect 140872 2984 140924 2990
rect 140872 2926 140924 2932
rect 141252 480 141280 3810
rect 146220 3806 146248 9454
rect 146312 9246 146340 12022
rect 147324 9450 147352 12022
rect 147312 9444 147364 9450
rect 147312 9386 147364 9392
rect 146300 9240 146352 9246
rect 146300 9182 146352 9188
rect 148336 8906 148364 12022
rect 149348 9382 149376 12022
rect 150452 9586 150480 12022
rect 150440 9580 150492 9586
rect 150440 9522 150492 9528
rect 151372 9518 151400 12022
rect 151912 9580 151964 9586
rect 151912 9522 151964 9528
rect 151360 9512 151412 9518
rect 151360 9454 151412 9460
rect 149336 9376 149388 9382
rect 149336 9318 149388 9324
rect 150440 9376 150492 9382
rect 150440 9318 150492 9324
rect 148968 9240 149020 9246
rect 148968 9182 149020 9188
rect 148324 8900 148376 8906
rect 148324 8842 148376 8848
rect 146944 8356 146996 8362
rect 146944 8298 146996 8304
rect 146208 3800 146260 3806
rect 146208 3742 146260 3748
rect 146956 3738 146984 8298
rect 147128 4072 147180 4078
rect 147128 4014 147180 4020
rect 146944 3732 146996 3738
rect 146944 3674 146996 3680
rect 142436 3528 142488 3534
rect 142436 3470 142488 3476
rect 142448 480 142476 3470
rect 143540 3460 143592 3466
rect 143540 3402 143592 3408
rect 143552 480 143580 3402
rect 145932 3324 145984 3330
rect 145932 3266 145984 3272
rect 144736 2984 144788 2990
rect 144736 2926 144788 2932
rect 144748 480 144776 2926
rect 145944 480 145972 3266
rect 147140 480 147168 4014
rect 148980 3874 149008 9182
rect 149704 8968 149756 8974
rect 149704 8910 149756 8916
rect 148968 3868 149020 3874
rect 148968 3810 149020 3816
rect 148324 3800 148376 3806
rect 148324 3742 148376 3748
rect 148336 480 148364 3742
rect 149520 3732 149572 3738
rect 149520 3674 149572 3680
rect 149532 480 149560 3674
rect 149716 3534 149744 8910
rect 149704 3528 149756 3534
rect 149704 3470 149756 3476
rect 150452 3466 150480 9318
rect 150716 9172 150768 9178
rect 150716 9114 150768 9120
rect 150624 3868 150676 3874
rect 150624 3810 150676 3816
rect 150440 3460 150492 3466
rect 150440 3402 150492 3408
rect 150636 480 150664 3810
rect 150728 2990 150756 9114
rect 151820 3460 151872 3466
rect 151820 3402 151872 3408
rect 150716 2984 150768 2990
rect 150716 2926 150768 2932
rect 151832 480 151860 3402
rect 151924 3330 151952 9522
rect 152384 8362 152412 12022
rect 153200 9444 153252 9450
rect 153200 9386 153252 9392
rect 152372 8356 152424 8362
rect 152372 8298 152424 8304
rect 153212 4078 153240 9386
rect 153396 9246 153424 12022
rect 153384 9240 153436 9246
rect 153384 9182 153436 9188
rect 154592 8974 154620 12022
rect 155420 9382 155448 12022
rect 155408 9376 155460 9382
rect 155408 9318 155460 9324
rect 156432 9178 156460 12022
rect 157444 9586 157472 12022
rect 157432 9580 157484 9586
rect 157432 9522 157484 9528
rect 157248 9512 157300 9518
rect 157248 9454 157300 9460
rect 156420 9172 156472 9178
rect 156420 9114 156472 9120
rect 155316 9104 155368 9110
rect 155316 9046 155368 9052
rect 154580 8968 154632 8974
rect 154580 8910 154632 8916
rect 153200 4072 153252 4078
rect 153200 4014 153252 4020
rect 155328 3806 155356 9046
rect 155316 3800 155368 3806
rect 155316 3742 155368 3748
rect 157260 3738 157288 9454
rect 158732 9450 158760 12022
rect 158720 9444 158772 9450
rect 158720 9386 158772 9392
rect 158996 9308 159048 9314
rect 158996 9250 159048 9256
rect 157708 9240 157760 9246
rect 157708 9182 157760 9188
rect 157720 3874 157748 9182
rect 158812 8356 158864 8362
rect 158812 8298 158864 8304
rect 157708 3868 157760 3874
rect 157708 3810 157760 3816
rect 157248 3732 157300 3738
rect 157248 3674 157300 3680
rect 157800 3732 157852 3738
rect 157800 3674 157852 3680
rect 154212 3664 154264 3670
rect 154212 3606 154264 3612
rect 153016 3528 153068 3534
rect 153016 3470 153068 3476
rect 151912 3324 151964 3330
rect 151912 3266 151964 3272
rect 153028 480 153056 3470
rect 154224 480 154252 3606
rect 156604 3596 156656 3602
rect 156604 3538 156656 3544
rect 155408 3324 155460 3330
rect 155408 3266 155460 3272
rect 155420 480 155448 3266
rect 156616 480 156644 3538
rect 157812 480 157840 3674
rect 158824 3466 158852 8298
rect 158904 3800 158956 3806
rect 158904 3742 158956 3748
rect 158812 3460 158864 3466
rect 158812 3402 158864 3408
rect 158916 480 158944 3742
rect 159008 3534 159036 9250
rect 159468 9110 159496 12022
rect 160480 9518 160508 12022
rect 160468 9512 160520 9518
rect 160468 9454 160520 9460
rect 161676 9246 161704 12022
rect 161664 9240 161716 9246
rect 161664 9182 161716 9188
rect 159456 9104 159508 9110
rect 159456 9046 159508 9052
rect 160100 9036 160152 9042
rect 160100 8978 160152 8984
rect 160112 3670 160140 8978
rect 161572 8764 161624 8770
rect 161572 8706 161624 8712
rect 161296 3868 161348 3874
rect 161296 3810 161348 3816
rect 160100 3664 160152 3670
rect 160100 3606 160152 3612
rect 158996 3528 159048 3534
rect 158996 3470 159048 3476
rect 160100 3460 160152 3466
rect 160100 3402 160152 3408
rect 160112 480 160140 3402
rect 161308 480 161336 3810
rect 161584 3330 161612 8706
rect 162504 8362 162532 12022
rect 163516 9314 163544 12022
rect 163504 9308 163556 9314
rect 163504 9250 163556 9256
rect 164528 9042 164556 12022
rect 165344 9444 165396 9450
rect 165344 9386 165396 9392
rect 164516 9036 164568 9042
rect 164516 8978 164568 8984
rect 162860 8900 162912 8906
rect 162860 8842 162912 8848
rect 162492 8356 162544 8362
rect 162492 8298 162544 8304
rect 162872 3602 162900 8842
rect 164884 4140 164936 4146
rect 164884 4082 164936 4088
rect 162860 3596 162912 3602
rect 162860 3538 162912 3544
rect 163688 3392 163740 3398
rect 163688 3334 163740 3340
rect 161572 3324 161624 3330
rect 161572 3266 161624 3272
rect 162492 2916 162544 2922
rect 162492 2858 162544 2864
rect 162504 480 162532 2858
rect 163700 480 163728 3334
rect 164896 480 164924 4082
rect 165356 3738 165384 9386
rect 165632 8770 165660 12022
rect 165988 9580 166040 9586
rect 165988 9522 166040 9528
rect 165620 8764 165672 8770
rect 165620 8706 165672 8712
rect 166000 3806 166028 9522
rect 166552 8906 166580 12022
rect 167276 9512 167328 9518
rect 167276 9454 167328 9460
rect 167092 9376 167144 9382
rect 167092 9318 167144 9324
rect 166540 8900 166592 8906
rect 166540 8842 166592 8848
rect 166080 4004 166132 4010
rect 166080 3946 166132 3952
rect 165988 3800 166040 3806
rect 165988 3742 166040 3748
rect 165344 3732 165396 3738
rect 165344 3674 165396 3680
rect 166092 480 166120 3946
rect 167104 3874 167132 9318
rect 167092 3868 167144 3874
rect 167092 3810 167144 3816
rect 167184 3800 167236 3806
rect 167184 3742 167236 3748
rect 167196 480 167224 3742
rect 167288 3466 167316 9454
rect 167564 9450 167592 12022
rect 168576 9586 168604 12022
rect 168564 9580 168616 9586
rect 168564 9522 168616 9528
rect 169772 9518 169800 12022
rect 169760 9512 169812 9518
rect 169760 9454 169812 9460
rect 167552 9444 167604 9450
rect 167552 9386 167604 9392
rect 170600 9382 170628 12022
rect 171232 9512 171284 9518
rect 171232 9454 171284 9460
rect 170588 9376 170640 9382
rect 170588 9318 170640 9324
rect 169944 9308 169996 9314
rect 169944 9250 169996 9256
rect 168472 8424 168524 8430
rect 168472 8366 168524 8372
rect 168380 3868 168432 3874
rect 168380 3810 168432 3816
rect 167276 3460 167328 3466
rect 167276 3402 167328 3408
rect 168392 480 168420 3810
rect 168484 2922 168512 8366
rect 169576 3460 169628 3466
rect 169576 3402 169628 3408
rect 168472 2916 168524 2922
rect 168472 2858 168524 2864
rect 169588 480 169616 3402
rect 169956 3398 169984 9250
rect 171244 4146 171272 9454
rect 171612 8430 171640 12022
rect 172624 9314 172652 12022
rect 173912 9518 173940 12022
rect 173900 9512 173952 9518
rect 173900 9454 173952 9460
rect 172612 9308 172664 9314
rect 172612 9250 172664 9256
rect 174648 8770 174676 12022
rect 175280 9512 175332 9518
rect 175280 9454 175332 9460
rect 175188 9444 175240 9450
rect 175188 9386 175240 9392
rect 172520 8764 172572 8770
rect 172520 8706 172572 8712
rect 174636 8764 174688 8770
rect 174636 8706 174688 8712
rect 171600 8424 171652 8430
rect 171600 8366 171652 8372
rect 171232 4140 171284 4146
rect 171232 4082 171284 4088
rect 172532 4010 172560 8706
rect 172520 4004 172572 4010
rect 172520 3946 172572 3952
rect 175200 3806 175228 9386
rect 175188 3800 175240 3806
rect 175188 3742 175240 3748
rect 170772 3664 170824 3670
rect 170772 3606 170824 3612
rect 169944 3392 169996 3398
rect 169944 3334 169996 3340
rect 170784 480 170812 3606
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 171968 2984 172020 2990
rect 171968 2926 172020 2932
rect 171980 480 172008 2926
rect 173176 480 173204 3470
rect 175292 3466 175320 9454
rect 175660 9450 175688 12022
rect 175648 9444 175700 9450
rect 175648 9386 175700 9392
rect 176672 8378 176700 12022
rect 177684 9518 177712 12022
rect 177672 9512 177724 9518
rect 177672 9454 177724 9460
rect 178696 9042 178724 12022
rect 179432 9466 179460 12022
rect 180812 9674 180840 12022
rect 179340 9438 179460 9466
rect 180720 9646 180840 9674
rect 177948 9036 178000 9042
rect 177948 8978 178000 8984
rect 178684 9036 178736 9042
rect 178684 8978 178736 8984
rect 176580 8350 176700 8378
rect 176580 3874 176608 8350
rect 176568 3868 176620 3874
rect 176568 3810 176620 3816
rect 176660 3868 176712 3874
rect 176660 3810 176712 3816
rect 175280 3460 175332 3466
rect 175280 3402 175332 3408
rect 174268 3324 174320 3330
rect 174268 3266 174320 3272
rect 174280 480 174308 3266
rect 175464 3188 175516 3194
rect 175464 3130 175516 3136
rect 175476 480 175504 3130
rect 176672 480 176700 3810
rect 177960 3670 177988 8978
rect 179052 3936 179104 3942
rect 179052 3878 179104 3884
rect 177948 3664 178000 3670
rect 177948 3606 178000 3612
rect 177856 3460 177908 3466
rect 177856 3402 177908 3408
rect 177868 480 177896 3402
rect 179064 480 179092 3878
rect 179340 2990 179368 9438
rect 180248 3596 180300 3602
rect 180248 3538 180300 3544
rect 179328 2984 179380 2990
rect 179328 2926 179380 2932
rect 180260 480 180288 3538
rect 180720 3534 180748 9646
rect 181272 6914 181300 12022
rect 180904 6886 181300 6914
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 180904 3330 180932 6886
rect 181444 3528 181496 3534
rect 181444 3470 181496 3476
rect 180892 3324 180944 3330
rect 180892 3266 180944 3272
rect 181456 480 181484 3470
rect 182192 3194 182220 12022
rect 183572 3874 183600 12022
rect 184952 9466 184980 12022
rect 184860 9438 184980 9466
rect 183560 3868 183612 3874
rect 183560 3810 183612 3816
rect 184860 3466 184888 9438
rect 185228 6914 185256 12022
rect 185136 6886 185256 6914
rect 184940 4004 184992 4010
rect 184940 3946 184992 3952
rect 184848 3460 184900 3466
rect 184848 3402 184900 3408
rect 182548 3324 182600 3330
rect 182548 3266 182600 3272
rect 182180 3188 182232 3194
rect 182180 3130 182232 3136
rect 182560 480 182588 3266
rect 183744 3188 183796 3194
rect 183744 3130 183796 3136
rect 183756 480 183784 3130
rect 184952 480 184980 3946
rect 185136 3942 185164 6886
rect 185124 3936 185176 3942
rect 185124 3878 185176 3884
rect 186332 3602 186360 12022
rect 186320 3596 186372 3602
rect 186320 3538 186372 3544
rect 187712 3534 187740 12022
rect 187700 3528 187752 3534
rect 187700 3470 187752 3476
rect 188528 3528 188580 3534
rect 188528 3470 188580 3476
rect 187332 3052 187384 3058
rect 187332 2994 187384 3000
rect 186136 2916 186188 2922
rect 186136 2858 186188 2864
rect 186148 480 186176 2858
rect 187344 480 187372 2994
rect 188540 480 188568 3470
rect 189092 3330 189120 12022
rect 189368 6914 189396 12022
rect 189184 6886 189396 6914
rect 189080 3324 189132 3330
rect 189080 3266 189132 3272
rect 189184 3194 189212 6886
rect 190472 4010 190500 12022
rect 190460 4004 190512 4010
rect 190460 3946 190512 3952
rect 189724 3732 189776 3738
rect 189724 3674 189776 3680
rect 189172 3188 189224 3194
rect 189172 3130 189224 3136
rect 189736 480 189764 3674
rect 190828 3460 190880 3466
rect 190828 3402 190880 3408
rect 190840 480 190868 3402
rect 191852 2922 191880 12022
rect 192312 6914 192340 12022
rect 193508 6914 193536 12022
rect 191944 6886 192340 6914
rect 193232 6886 193536 6914
rect 191944 3058 191972 6886
rect 193232 3534 193260 6886
rect 194612 3738 194640 12022
rect 195612 4004 195664 4010
rect 195612 3946 195664 3952
rect 194600 3732 194652 3738
rect 194600 3674 194652 3680
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 194416 3528 194468 3534
rect 194416 3470 194468 3476
rect 192024 3324 192076 3330
rect 192024 3266 192076 3272
rect 191932 3052 191984 3058
rect 191932 2994 191984 3000
rect 191840 2916 191892 2922
rect 191840 2858 191892 2864
rect 192036 480 192064 3266
rect 193220 3256 193272 3262
rect 193220 3198 193272 3204
rect 193232 480 193260 3198
rect 194428 480 194456 3470
rect 195624 480 195652 3946
rect 195992 3466 196020 12022
rect 196360 6914 196388 12022
rect 196084 6886 196388 6914
rect 195980 3460 196032 3466
rect 195980 3402 196032 3408
rect 196084 3330 196112 6886
rect 196808 3800 196860 3806
rect 196808 3742 196860 3748
rect 196072 3324 196124 3330
rect 196072 3266 196124 3272
rect 196820 480 196848 3742
rect 197372 3262 197400 12022
rect 197912 4140 197964 4146
rect 197912 4082 197964 4088
rect 197360 3256 197412 3262
rect 197360 3198 197412 3204
rect 197924 480 197952 4082
rect 198752 3534 198780 12022
rect 200120 9512 200172 9518
rect 200120 9454 200172 9460
rect 200132 3806 200160 9454
rect 200224 4010 200252 12022
rect 200960 9518 200988 12022
rect 200948 9512 201000 9518
rect 200948 9454 201000 9460
rect 201500 9512 201552 9518
rect 201500 9454 201552 9460
rect 200212 4004 200264 4010
rect 200212 3946 200264 3952
rect 200120 3800 200172 3806
rect 200120 3742 200172 3748
rect 199108 3732 199160 3738
rect 199108 3674 199160 3680
rect 198740 3528 198792 3534
rect 198740 3470 198792 3476
rect 199120 480 199148 3674
rect 200304 3528 200356 3534
rect 200304 3470 200356 3476
rect 200316 480 200344 3470
rect 201512 480 201540 9454
rect 201604 4146 201632 12022
rect 201592 4140 201644 4146
rect 201592 4082 201644 4088
rect 202892 3738 202920 12022
rect 204318 11778 204346 12036
rect 205008 12022 205344 12050
rect 205744 12022 206356 12050
rect 207124 12022 207368 12050
rect 208044 12022 208380 12050
rect 209056 12022 209392 12050
rect 210068 12022 210404 12050
rect 211172 12022 211416 12050
rect 212092 12022 212428 12050
rect 213104 12022 213440 12050
rect 214116 12022 214452 12050
rect 215312 12022 215464 12050
rect 216140 12022 216476 12050
rect 217152 12022 217488 12050
rect 218164 12022 218500 12050
rect 204318 11750 204392 11778
rect 202880 3732 202932 3738
rect 202880 3674 202932 3680
rect 204364 3534 204392 11750
rect 205008 9518 205036 12022
rect 204996 9512 205048 9518
rect 204996 9454 205048 9460
rect 205088 8764 205140 8770
rect 205088 8706 205140 8712
rect 204352 3528 204404 3534
rect 204352 3470 204404 3476
rect 202696 3324 202748 3330
rect 202696 3266 202748 3272
rect 202708 480 202736 3266
rect 203892 3256 203944 3262
rect 203892 3198 203944 3204
rect 203904 480 203932 3198
rect 205100 480 205128 8706
rect 205744 3330 205772 12022
rect 206192 9512 206244 9518
rect 206192 9454 206244 9460
rect 205732 3324 205784 3330
rect 205732 3266 205784 3272
rect 206204 480 206232 9454
rect 207124 3262 207152 12022
rect 208044 8770 208072 12022
rect 209056 9518 209084 12022
rect 209044 9512 209096 9518
rect 209044 9454 209096 9460
rect 209780 9036 209832 9042
rect 209780 8978 209832 8984
rect 208032 8764 208084 8770
rect 208032 8706 208084 8712
rect 207388 8492 207440 8498
rect 207388 8434 207440 8440
rect 207112 3256 207164 3262
rect 207112 3198 207164 3204
rect 207400 480 207428 8434
rect 208584 8424 208636 8430
rect 208584 8366 208636 8372
rect 208596 480 208624 8366
rect 209792 480 209820 8978
rect 210068 8498 210096 12022
rect 210976 9512 211028 9518
rect 210976 9454 211028 9460
rect 210056 8492 210108 8498
rect 210056 8434 210108 8440
rect 210988 480 211016 9454
rect 211172 8430 211200 12022
rect 212092 9042 212120 12022
rect 213104 9518 213132 12022
rect 213092 9512 213144 9518
rect 213092 9454 213144 9460
rect 213368 9512 213420 9518
rect 213368 9454 213420 9460
rect 212080 9036 212132 9042
rect 212080 8978 212132 8984
rect 212172 8560 212224 8566
rect 212172 8502 212224 8508
rect 211160 8424 211212 8430
rect 211160 8366 211212 8372
rect 212184 480 212212 8502
rect 213380 480 213408 9454
rect 214116 8566 214144 12022
rect 215312 9518 215340 12022
rect 215300 9512 215352 9518
rect 215300 9454 215352 9460
rect 215668 9512 215720 9518
rect 215668 9454 215720 9460
rect 214472 8900 214524 8906
rect 214472 8842 214524 8848
rect 214104 8560 214156 8566
rect 214104 8502 214156 8508
rect 214484 480 214512 8842
rect 215680 480 215708 9454
rect 216140 8906 216168 12022
rect 217152 9518 217180 12022
rect 217140 9512 217192 9518
rect 217140 9454 217192 9460
rect 218164 9314 218192 12022
rect 219498 11778 219526 12036
rect 220188 12022 220524 12050
rect 221200 12022 221536 12050
rect 222212 12022 222548 12050
rect 222764 12022 223560 12050
rect 223684 12022 224572 12050
rect 225156 12022 225584 12050
rect 226352 12022 226596 12050
rect 227548 12022 227608 12050
rect 228284 12022 228620 12050
rect 229388 12022 229632 12050
rect 230644 12022 231072 12050
rect 231656 12022 231808 12050
rect 232668 12022 233004 12050
rect 233680 12022 234016 12050
rect 219498 11750 219572 11778
rect 219268 9654 219480 9674
rect 219268 9648 219492 9654
rect 219268 9646 219440 9648
rect 216864 9308 216916 9314
rect 216864 9250 216916 9256
rect 218152 9308 218204 9314
rect 218152 9250 218204 9256
rect 216128 8900 216180 8906
rect 216128 8842 216180 8848
rect 216876 480 216904 9250
rect 218060 8356 218112 8362
rect 218060 8298 218112 8304
rect 218072 480 218100 8298
rect 219268 480 219296 9646
rect 219440 9590 219492 9596
rect 219544 8362 219572 11750
rect 220188 9654 220216 12022
rect 220176 9648 220228 9654
rect 220176 9590 220228 9596
rect 221200 8770 221228 12022
rect 222212 9450 222240 12022
rect 221556 9444 221608 9450
rect 221556 9386 221608 9392
rect 222200 9444 222252 9450
rect 222200 9386 222252 9392
rect 220452 8764 220504 8770
rect 220452 8706 220504 8712
rect 221188 8764 221240 8770
rect 221188 8706 221240 8712
rect 219532 8356 219584 8362
rect 219532 8298 219584 8304
rect 220464 480 220492 8706
rect 221568 480 221596 9386
rect 222764 480 222792 12022
rect 223684 6914 223712 12022
rect 223592 6886 223712 6914
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223592 354 223620 6886
rect 225156 480 225184 12022
rect 226352 480 226380 12022
rect 227548 480 227576 12022
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 12022
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 12022
rect 231044 480 231072 12022
rect 231780 9518 231808 12022
rect 232976 9518 233004 12022
rect 233988 9518 234016 12022
rect 234632 12022 234692 12050
rect 235704 12022 235948 12050
rect 236716 12022 236960 12050
rect 237728 12022 238064 12050
rect 231768 9512 231820 9518
rect 231768 9454 231820 9460
rect 232228 9512 232280 9518
rect 232228 9454 232280 9460
rect 232964 9512 233016 9518
rect 232964 9454 233016 9460
rect 233424 9512 233476 9518
rect 233424 9454 233476 9460
rect 233976 9512 234028 9518
rect 233976 9454 234028 9460
rect 232240 480 232268 9454
rect 233436 480 233464 9454
rect 234632 3602 234660 12022
rect 235920 9518 235948 12022
rect 234712 9512 234764 9518
rect 234712 9454 234764 9460
rect 235908 9512 235960 9518
rect 235908 9454 235960 9460
rect 234620 3596 234672 3602
rect 234620 3538 234672 3544
rect 234724 3482 234752 9454
rect 236932 9450 236960 12022
rect 237012 9512 237064 9518
rect 237012 9454 237064 9460
rect 236920 9444 236972 9450
rect 236920 9386 236972 9392
rect 235816 3596 235868 3602
rect 235816 3538 235868 3544
rect 234632 3454 234752 3482
rect 234632 480 234660 3454
rect 235828 480 235856 3538
rect 237024 480 237052 9454
rect 238036 8362 238064 12022
rect 238680 12022 238740 12050
rect 239752 12022 240088 12050
rect 240764 12022 241100 12050
rect 241776 12022 242112 12050
rect 238116 9444 238168 9450
rect 238116 9386 238168 9392
rect 238024 8356 238076 8362
rect 238024 8298 238076 8304
rect 238128 480 238156 9386
rect 238680 8498 238708 12022
rect 240060 9466 240088 12022
rect 240060 9438 240272 9466
rect 238668 8492 238720 8498
rect 238668 8434 238720 8440
rect 240048 8492 240100 8498
rect 240048 8434 240100 8440
rect 239312 8356 239364 8362
rect 239312 8298 239364 8304
rect 239324 480 239352 8298
rect 240060 2802 240088 8434
rect 240244 3534 240272 9438
rect 241072 9382 241100 12022
rect 241060 9376 241112 9382
rect 241060 9318 241112 9324
rect 242084 8634 242112 12022
rect 242728 12022 242788 12050
rect 243800 12022 244136 12050
rect 244812 12022 245148 12050
rect 245824 12022 246160 12050
rect 246836 12022 246988 12050
rect 247848 12022 248184 12050
rect 248860 12022 249196 12050
rect 249872 12022 250208 12050
rect 250884 12022 251128 12050
rect 251896 12022 252232 12050
rect 252908 12022 253244 12050
rect 242728 8906 242756 12022
rect 242808 9376 242860 9382
rect 242808 9318 242860 9324
rect 242716 8900 242768 8906
rect 242716 8842 242768 8848
rect 242072 8628 242124 8634
rect 242072 8570 242124 8576
rect 240232 3528 240284 3534
rect 240232 3470 240284 3476
rect 241704 3528 241756 3534
rect 241704 3470 241756 3476
rect 242820 3482 242848 9318
rect 243268 8900 243320 8906
rect 243268 8842 243320 8848
rect 240060 2774 240180 2802
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 354 240180 2774
rect 241716 480 241744 3470
rect 242820 3454 242940 3482
rect 242912 480 242940 3454
rect 243280 3058 243308 8842
rect 244108 8770 244136 12022
rect 245120 9518 245148 12022
rect 245108 9512 245160 9518
rect 245108 9454 245160 9460
rect 245844 9512 245896 9518
rect 245844 9454 245896 9460
rect 244096 8764 244148 8770
rect 244096 8706 244148 8712
rect 244648 8764 244700 8770
rect 244648 8706 244700 8712
rect 244096 8628 244148 8634
rect 244096 8570 244148 8576
rect 243268 3052 243320 3058
rect 243268 2994 243320 3000
rect 244108 480 244136 8570
rect 244660 3534 244688 8706
rect 244648 3528 244700 3534
rect 244648 3470 244700 3476
rect 245856 3058 245884 9454
rect 246132 9178 246160 12022
rect 246960 9450 246988 12022
rect 246948 9444 247000 9450
rect 246948 9386 247000 9392
rect 247868 9444 247920 9450
rect 247868 9386 247920 9392
rect 246120 9172 246172 9178
rect 246120 9114 246172 9120
rect 247880 4146 247908 9386
rect 248156 8702 248184 12022
rect 249168 9314 249196 12022
rect 249156 9308 249208 9314
rect 249156 9250 249208 9256
rect 249800 9308 249852 9314
rect 249800 9250 249852 9256
rect 248328 9172 248380 9178
rect 248328 9114 248380 9120
rect 248144 8696 248196 8702
rect 248144 8638 248196 8644
rect 247868 4140 247920 4146
rect 247868 4082 247920 4088
rect 246396 3528 246448 3534
rect 246396 3470 246448 3476
rect 245200 3052 245252 3058
rect 245200 2994 245252 3000
rect 245844 3052 245896 3058
rect 245844 2994 245896 3000
rect 245212 480 245240 2994
rect 246408 480 246436 3470
rect 247592 3052 247644 3058
rect 247592 2994 247644 3000
rect 247604 480 247632 2994
rect 248340 2802 248368 9114
rect 248512 8696 248564 8702
rect 248512 8638 248564 8644
rect 248524 3330 248552 8638
rect 249812 3534 249840 9250
rect 250180 8634 250208 12022
rect 251100 9518 251128 12022
rect 251088 9512 251140 9518
rect 251088 9454 251140 9460
rect 252204 9450 252232 12022
rect 252284 9512 252336 9518
rect 252284 9454 252336 9460
rect 252192 9444 252244 9450
rect 252192 9386 252244 9392
rect 250168 8628 250220 8634
rect 250168 8570 250220 8576
rect 249984 4140 250036 4146
rect 249984 4082 250036 4088
rect 249800 3528 249852 3534
rect 249800 3470 249852 3476
rect 248512 3324 248564 3330
rect 248512 3266 248564 3272
rect 248340 2774 248460 2802
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 2774
rect 249996 480 250024 4082
rect 251180 3324 251232 3330
rect 251180 3266 251232 3272
rect 251192 480 251220 3266
rect 252296 3058 252324 9454
rect 253216 8770 253244 12022
rect 253860 12022 253920 12050
rect 254932 12022 255176 12050
rect 255944 12022 256280 12050
rect 256956 12022 257292 12050
rect 253860 9518 253888 12022
rect 253848 9512 253900 9518
rect 253848 9454 253900 9460
rect 253480 9444 253532 9450
rect 253480 9386 253532 9392
rect 253204 8764 253256 8770
rect 253204 8706 253256 8712
rect 252468 8628 252520 8634
rect 252468 8570 252520 8576
rect 252480 3534 252508 8570
rect 253492 3670 253520 9386
rect 255148 8906 255176 12022
rect 256252 9518 256280 12022
rect 255228 9512 255280 9518
rect 255228 9454 255280 9460
rect 256240 9512 256292 9518
rect 256240 9454 256292 9460
rect 255136 8900 255188 8906
rect 255136 8842 255188 8848
rect 254768 8764 254820 8770
rect 254768 8706 254820 8712
rect 253480 3664 253532 3670
rect 253480 3606 253532 3612
rect 252376 3528 252428 3534
rect 252376 3470 252428 3476
rect 252468 3528 252520 3534
rect 252468 3470 252520 3476
rect 253480 3528 253532 3534
rect 253480 3470 253532 3476
rect 252284 3052 252336 3058
rect 252284 2994 252336 3000
rect 252388 480 252416 3470
rect 253492 480 253520 3470
rect 254780 3194 254808 8706
rect 255240 4010 255268 9454
rect 256608 8900 256660 8906
rect 256608 8842 256660 8848
rect 255228 4004 255280 4010
rect 255228 3946 255280 3952
rect 255872 3664 255924 3670
rect 255872 3606 255924 3612
rect 254768 3188 254820 3194
rect 254768 3130 254820 3136
rect 254676 3052 254728 3058
rect 254676 2994 254728 3000
rect 254688 480 254716 2994
rect 255884 480 255912 3606
rect 256620 3466 256648 8842
rect 257264 8566 257292 12022
rect 257954 11778 257982 12036
rect 258980 12022 259408 12050
rect 259992 12022 260328 12050
rect 261004 12022 261340 12050
rect 262016 12022 262168 12050
rect 263028 12022 263364 12050
rect 264040 12022 264376 12050
rect 265052 12022 265388 12050
rect 266064 12022 266308 12050
rect 267076 12022 267412 12050
rect 268088 12022 268424 12050
rect 257954 11750 258028 11778
rect 257896 9512 257948 9518
rect 257896 9454 257948 9460
rect 257252 8560 257304 8566
rect 257252 8502 257304 8508
rect 257908 3874 257936 9454
rect 258000 9246 258028 11750
rect 259380 9466 259408 12022
rect 259380 9438 259500 9466
rect 257988 9240 258040 9246
rect 257988 9182 258040 9188
rect 258172 9240 258224 9246
rect 258172 9182 258224 9188
rect 258080 8560 258132 8566
rect 258080 8502 258132 8508
rect 257896 3868 257948 3874
rect 257896 3810 257948 3816
rect 258092 3534 258120 8502
rect 258184 3602 258212 9182
rect 258264 4004 258316 4010
rect 258264 3946 258316 3952
rect 258172 3596 258224 3602
rect 258172 3538 258224 3544
rect 258080 3528 258132 3534
rect 258080 3470 258132 3476
rect 256608 3460 256660 3466
rect 256608 3402 256660 3408
rect 257068 3188 257120 3194
rect 257068 3130 257120 3136
rect 257080 480 257108 3130
rect 258276 480 258304 3946
rect 259472 3670 259500 9438
rect 260300 9382 260328 12022
rect 261312 9586 261340 12022
rect 261300 9580 261352 9586
rect 261300 9522 261352 9528
rect 262140 9518 262168 12022
rect 262128 9512 262180 9518
rect 262128 9454 262180 9460
rect 263336 9450 263364 12022
rect 263508 9580 263560 9586
rect 263508 9522 263560 9528
rect 263416 9512 263468 9518
rect 263416 9454 263468 9460
rect 263324 9444 263376 9450
rect 263324 9386 263376 9392
rect 260288 9376 260340 9382
rect 260288 9318 260340 9324
rect 262128 9376 262180 9382
rect 262128 9318 262180 9324
rect 260656 3868 260708 3874
rect 260656 3810 260708 3816
rect 259460 3664 259512 3670
rect 259460 3606 259512 3612
rect 259460 3460 259512 3466
rect 259460 3402 259512 3408
rect 259472 480 259500 3402
rect 260668 480 260696 3810
rect 261760 3528 261812 3534
rect 261760 3470 261812 3476
rect 261772 480 261800 3470
rect 262140 3262 262168 9318
rect 262956 3596 263008 3602
rect 262956 3538 263008 3544
rect 262128 3256 262180 3262
rect 262128 3198 262180 3204
rect 262968 480 262996 3538
rect 263428 3398 263456 9454
rect 263520 3534 263548 9522
rect 264348 8770 264376 12022
rect 265360 9518 265388 12022
rect 265348 9512 265400 9518
rect 265348 9454 265400 9460
rect 264888 9444 264940 9450
rect 264888 9386 264940 9392
rect 264336 8764 264388 8770
rect 264336 8706 264388 8712
rect 264900 3874 264928 9386
rect 266280 8906 266308 12022
rect 266268 8900 266320 8906
rect 266268 8842 266320 8848
rect 266728 8900 266780 8906
rect 266728 8842 266780 8848
rect 266268 8764 266320 8770
rect 266268 8706 266320 8712
rect 264888 3868 264940 3874
rect 264888 3810 264940 3816
rect 264152 3664 264204 3670
rect 264152 3606 264204 3612
rect 263508 3528 263560 3534
rect 263508 3470 263560 3476
rect 263416 3392 263468 3398
rect 263416 3334 263468 3340
rect 264164 480 264192 3606
rect 266280 3330 266308 8706
rect 266740 3602 266768 8842
rect 267384 8702 267412 12022
rect 267648 9512 267700 9518
rect 267648 9454 267700 9460
rect 267372 8696 267424 8702
rect 267372 8638 267424 8644
rect 267660 3806 267688 9454
rect 268396 9042 268424 12022
rect 269040 12022 269100 12050
rect 270112 12022 270448 12050
rect 271124 12022 271460 12050
rect 272136 12022 272472 12050
rect 269040 9466 269068 12022
rect 269040 9438 269252 9466
rect 268384 9036 268436 9042
rect 268384 8978 268436 8984
rect 269120 9036 269172 9042
rect 269120 8978 269172 8984
rect 267740 8696 267792 8702
rect 267740 8638 267792 8644
rect 267648 3800 267700 3806
rect 267648 3742 267700 3748
rect 267752 3670 267780 8638
rect 268844 3868 268896 3874
rect 268844 3810 268896 3816
rect 267740 3664 267792 3670
rect 267740 3606 267792 3612
rect 266728 3596 266780 3602
rect 266728 3538 266780 3544
rect 266544 3528 266596 3534
rect 266544 3470 266596 3476
rect 266268 3324 266320 3330
rect 266268 3266 266320 3272
rect 265348 3256 265400 3262
rect 265348 3198 265400 3204
rect 265360 480 265388 3198
rect 266556 480 266584 3470
rect 267740 3392 267792 3398
rect 267740 3334 267792 3340
rect 267752 480 267780 3334
rect 268856 480 268884 3810
rect 269132 3534 269160 8978
rect 269120 3528 269172 3534
rect 269120 3470 269172 3476
rect 269224 2990 269252 9438
rect 270420 8770 270448 12022
rect 271432 9382 271460 12022
rect 271420 9376 271472 9382
rect 271420 9318 271472 9324
rect 272444 9314 272472 12022
rect 273088 12022 273148 12050
rect 274160 12022 274496 12050
rect 275172 12022 275508 12050
rect 276184 12022 276520 12050
rect 277196 12022 277348 12050
rect 278208 12022 278728 12050
rect 279220 12022 279556 12050
rect 280232 12022 280568 12050
rect 281244 12022 281488 12050
rect 282256 12022 282592 12050
rect 283268 12022 283604 12050
rect 273088 9518 273116 12022
rect 273076 9512 273128 9518
rect 273076 9454 273128 9460
rect 274468 9450 274496 12022
rect 275480 9518 275508 12022
rect 274548 9512 274600 9518
rect 274548 9454 274600 9460
rect 275468 9512 275520 9518
rect 275468 9454 275520 9460
rect 274456 9444 274508 9450
rect 274456 9386 274508 9392
rect 273168 9376 273220 9382
rect 273168 9318 273220 9324
rect 272432 9308 272484 9314
rect 272432 9250 272484 9256
rect 270408 8764 270460 8770
rect 270408 8706 270460 8712
rect 271788 8764 271840 8770
rect 271788 8706 271840 8712
rect 271236 3800 271288 3806
rect 271236 3742 271288 3748
rect 270040 3324 270092 3330
rect 270040 3266 270092 3272
rect 269212 2984 269264 2990
rect 269212 2926 269264 2932
rect 270052 480 270080 3266
rect 271248 480 271276 3742
rect 271800 3330 271828 8706
rect 273180 4010 273208 9318
rect 274456 9308 274508 9314
rect 274456 9250 274508 9256
rect 274468 4146 274496 9250
rect 274456 4140 274508 4146
rect 274456 4082 274508 4088
rect 273168 4004 273220 4010
rect 273168 3946 273220 3952
rect 274560 3806 274588 9454
rect 275836 9444 275888 9450
rect 275836 9386 275888 9392
rect 274548 3800 274600 3806
rect 274548 3742 274600 3748
rect 273628 3664 273680 3670
rect 273628 3606 273680 3612
rect 272432 3596 272484 3602
rect 272432 3538 272484 3544
rect 271788 3324 271840 3330
rect 271788 3266 271840 3272
rect 272444 480 272472 3538
rect 273640 480 273668 3606
rect 275848 3534 275876 9386
rect 276492 8566 276520 12022
rect 276756 9512 276808 9518
rect 276756 9454 276808 9460
rect 276480 8560 276532 8566
rect 276480 8502 276532 8508
rect 274824 3528 274876 3534
rect 274824 3470 274876 3476
rect 275836 3528 275888 3534
rect 275836 3470 275888 3476
rect 274836 480 274864 3470
rect 276768 3466 276796 9454
rect 277320 9110 277348 12022
rect 278700 9466 278728 12022
rect 278700 9438 278820 9466
rect 277308 9104 277360 9110
rect 277308 9046 277360 9052
rect 277676 9104 277728 9110
rect 277676 9046 277728 9052
rect 277400 8560 277452 8566
rect 277400 8502 277452 8508
rect 276756 3460 276808 3466
rect 276756 3402 276808 3408
rect 277412 3398 277440 8502
rect 277400 3392 277452 3398
rect 277400 3334 277452 3340
rect 277124 3324 277176 3330
rect 277124 3266 277176 3272
rect 276020 2984 276072 2990
rect 276020 2926 276072 2932
rect 276032 480 276060 2926
rect 277136 480 277164 3266
rect 277688 3058 277716 9046
rect 278320 4004 278372 4010
rect 278320 3946 278372 3952
rect 277676 3052 277728 3058
rect 277676 2994 277728 3000
rect 278332 480 278360 3946
rect 278792 3670 278820 9438
rect 279528 8566 279556 12022
rect 280540 9518 280568 12022
rect 280528 9512 280580 9518
rect 280528 9454 280580 9460
rect 281460 8702 281488 12022
rect 282564 9178 282592 12022
rect 283576 9518 283604 12022
rect 284220 12022 284280 12050
rect 285292 12022 285628 12050
rect 286304 12022 286640 12050
rect 287316 12022 287652 12050
rect 282828 9512 282880 9518
rect 282828 9454 282880 9460
rect 283564 9512 283616 9518
rect 283564 9454 283616 9460
rect 282552 9172 282604 9178
rect 282552 9114 282604 9120
rect 281448 8696 281500 8702
rect 281448 8638 281500 8644
rect 282736 8696 282788 8702
rect 282736 8638 282788 8644
rect 279516 8560 279568 8566
rect 279516 8502 279568 8508
rect 281448 8560 281500 8566
rect 281448 8502 281500 8508
rect 281460 4146 281488 8502
rect 279516 4140 279568 4146
rect 279516 4082 279568 4088
rect 281448 4140 281500 4146
rect 281448 4082 281500 4088
rect 278780 3664 278832 3670
rect 278780 3606 278832 3612
rect 279528 480 279556 4082
rect 280712 3800 280764 3806
rect 280712 3742 280764 3748
rect 280724 480 280752 3742
rect 282748 3534 282776 8638
rect 282840 4078 282868 9454
rect 284220 9314 284248 12022
rect 285496 9512 285548 9518
rect 285496 9454 285548 9460
rect 284208 9308 284260 9314
rect 284208 9250 284260 9256
rect 284208 9172 284260 9178
rect 284208 9114 284260 9120
rect 282828 4072 282880 4078
rect 282828 4014 282880 4020
rect 284220 3874 284248 9114
rect 284208 3868 284260 3874
rect 284208 3810 284260 3816
rect 285508 3602 285536 9454
rect 285600 9450 285628 12022
rect 285588 9444 285640 9450
rect 285588 9386 285640 9392
rect 286140 9444 286192 9450
rect 286140 9386 286192 9392
rect 285588 9308 285640 9314
rect 285588 9250 285640 9256
rect 285600 3942 285628 9250
rect 285588 3936 285640 3942
rect 285588 3878 285640 3884
rect 286152 3738 286180 9386
rect 286612 8974 286640 12022
rect 287624 9518 287652 12022
rect 288314 11778 288342 12036
rect 289340 12022 289676 12050
rect 290352 12022 290688 12050
rect 291364 12022 291700 12050
rect 292376 12022 292528 12050
rect 293388 12022 293724 12050
rect 294400 12022 294736 12050
rect 295412 12022 295748 12050
rect 296424 12022 296576 12050
rect 297436 12022 298048 12050
rect 298448 12022 298784 12050
rect 288314 11750 288388 11778
rect 287612 9512 287664 9518
rect 287612 9454 287664 9460
rect 288360 9466 288388 11750
rect 288532 9512 288584 9518
rect 288360 9438 288480 9466
rect 288532 9454 288584 9460
rect 286600 8968 286652 8974
rect 286600 8910 286652 8916
rect 287336 8968 287388 8974
rect 287336 8910 287388 8916
rect 286140 3732 286192 3738
rect 286140 3674 286192 3680
rect 286600 3664 286652 3670
rect 286600 3606 286652 3612
rect 285496 3596 285548 3602
rect 285496 3538 285548 3544
rect 281908 3528 281960 3534
rect 281908 3470 281960 3476
rect 282736 3528 282788 3534
rect 282736 3470 282788 3476
rect 281920 480 281948 3470
rect 283104 3460 283156 3466
rect 283104 3402 283156 3408
rect 283116 480 283144 3402
rect 284300 3392 284352 3398
rect 284300 3334 284352 3340
rect 284312 480 284340 3334
rect 285404 3052 285456 3058
rect 285404 2994 285456 3000
rect 285416 480 285444 2994
rect 286612 480 286640 3606
rect 287348 3058 287376 8910
rect 287796 4140 287848 4146
rect 287796 4082 287848 4088
rect 287336 3052 287388 3058
rect 287336 2994 287388 3000
rect 287808 480 287836 4082
rect 288452 3670 288480 9438
rect 288440 3664 288492 3670
rect 288440 3606 288492 3612
rect 288544 3466 288572 9454
rect 289648 9178 289676 12022
rect 290660 9382 290688 12022
rect 290648 9376 290700 9382
rect 290648 9318 290700 9324
rect 289636 9172 289688 9178
rect 289636 9114 289688 9120
rect 290832 9172 290884 9178
rect 290832 9114 290884 9120
rect 288992 4072 289044 4078
rect 288992 4014 289044 4020
rect 288532 3460 288584 3466
rect 288532 3402 288584 3408
rect 289004 480 289032 4014
rect 290844 3534 290872 9114
rect 291672 9042 291700 12022
rect 292500 9518 292528 12022
rect 292488 9512 292540 9518
rect 292488 9454 292540 9460
rect 292488 9376 292540 9382
rect 292488 9318 292540 9324
rect 291660 9036 291712 9042
rect 291660 8978 291712 8984
rect 292500 3874 292528 9318
rect 293696 8634 293724 12022
rect 293868 9512 293920 9518
rect 293868 9454 293920 9460
rect 293776 9036 293828 9042
rect 293776 8978 293828 8984
rect 293684 8628 293736 8634
rect 293684 8570 293736 8576
rect 293684 3936 293736 3942
rect 293684 3878 293736 3884
rect 291384 3868 291436 3874
rect 291384 3810 291436 3816
rect 292488 3868 292540 3874
rect 292488 3810 292540 3816
rect 290188 3528 290240 3534
rect 290188 3470 290240 3476
rect 290832 3528 290884 3534
rect 290832 3470 290884 3476
rect 290200 480 290228 3470
rect 291396 480 291424 3810
rect 292580 3596 292632 3602
rect 292580 3538 292632 3544
rect 292592 480 292620 3538
rect 293696 480 293724 3878
rect 293788 3398 293816 8978
rect 293880 3602 293908 9454
rect 294708 9450 294736 12022
rect 294696 9444 294748 9450
rect 294696 9386 294748 9392
rect 295064 8628 295116 8634
rect 295064 8570 295116 8576
rect 295076 3738 295104 8570
rect 295720 8362 295748 12022
rect 295892 9444 295944 9450
rect 295892 9386 295944 9392
rect 295708 8356 295760 8362
rect 295708 8298 295760 8304
rect 295904 4010 295932 9386
rect 296548 8430 296576 12022
rect 298020 9466 298048 12022
rect 298020 9438 298140 9466
rect 296536 8424 296588 8430
rect 296536 8366 296588 8372
rect 297456 8424 297508 8430
rect 297456 8366 297508 8372
rect 296720 8356 296772 8362
rect 296720 8298 296772 8304
rect 296732 4078 296760 8298
rect 296720 4072 296772 4078
rect 296720 4014 296772 4020
rect 295892 4004 295944 4010
rect 295892 3946 295944 3952
rect 294880 3732 294932 3738
rect 294880 3674 294932 3680
rect 295064 3732 295116 3738
rect 295064 3674 295116 3680
rect 293868 3596 293920 3602
rect 293868 3538 293920 3544
rect 293776 3392 293828 3398
rect 293776 3334 293828 3340
rect 294892 480 294920 3674
rect 297468 3466 297496 8366
rect 298112 3806 298140 9438
rect 298756 9246 298784 12022
rect 299400 12022 299460 12050
rect 300472 12022 300808 12050
rect 301484 12022 301820 12050
rect 302496 12022 302832 12050
rect 299400 9314 299428 12022
rect 300780 9450 300808 12022
rect 301792 9518 301820 12022
rect 301780 9512 301832 9518
rect 301780 9454 301832 9460
rect 300768 9444 300820 9450
rect 300768 9386 300820 9392
rect 302148 9444 302200 9450
rect 302148 9386 302200 9392
rect 299388 9308 299440 9314
rect 299388 9250 299440 9256
rect 299940 9308 299992 9314
rect 299940 9250 299992 9256
rect 298744 9240 298796 9246
rect 298744 9182 298796 9188
rect 299952 3942 299980 9250
rect 300768 9240 300820 9246
rect 300768 9182 300820 9188
rect 300780 4146 300808 9182
rect 300768 4140 300820 4146
rect 300768 4082 300820 4088
rect 299940 3936 299992 3942
rect 299940 3878 299992 3884
rect 300768 3868 300820 3874
rect 300768 3810 300820 3816
rect 298100 3800 298152 3806
rect 298100 3742 298152 3748
rect 298468 3664 298520 3670
rect 298468 3606 298520 3612
rect 297272 3460 297324 3466
rect 297272 3402 297324 3408
rect 297456 3460 297508 3466
rect 297456 3402 297508 3408
rect 296076 3052 296128 3058
rect 296076 2994 296128 3000
rect 296088 480 296116 2994
rect 297284 480 297312 3402
rect 298480 480 298508 3606
rect 299664 3528 299716 3534
rect 299664 3470 299716 3476
rect 299676 480 299704 3470
rect 300780 480 300808 3810
rect 302160 3806 302188 9386
rect 302804 9042 302832 12022
rect 303448 12022 303508 12050
rect 304520 12022 304856 12050
rect 305532 12022 305868 12050
rect 306544 12022 306880 12050
rect 307556 12022 307708 12050
rect 308568 12022 308904 12050
rect 309580 12022 309916 12050
rect 310592 12022 310928 12050
rect 311604 12022 311848 12050
rect 312616 12022 312952 12050
rect 313628 12022 313964 12050
rect 303068 9512 303120 9518
rect 303068 9454 303120 9460
rect 302792 9036 302844 9042
rect 302792 8978 302844 8984
rect 302148 3800 302200 3806
rect 302148 3742 302200 3748
rect 303080 3670 303108 9454
rect 303448 8974 303476 12022
rect 304828 9450 304856 12022
rect 304816 9444 304868 9450
rect 304816 9386 304868 9392
rect 304908 9036 304960 9042
rect 304908 8978 304960 8984
rect 303436 8968 303488 8974
rect 303436 8910 303488 8916
rect 304356 3732 304408 3738
rect 304356 3674 304408 3680
rect 303068 3664 303120 3670
rect 303068 3606 303120 3612
rect 303160 3596 303212 3602
rect 303160 3538 303212 3544
rect 301964 3392 302016 3398
rect 301964 3334 302016 3340
rect 301976 480 302004 3334
rect 303172 480 303200 3538
rect 304368 480 304396 3674
rect 304920 3602 304948 8978
rect 305840 8430 305868 12022
rect 306852 9518 306880 12022
rect 307680 9586 307708 12022
rect 307668 9580 307720 9586
rect 307668 9522 307720 9528
rect 306840 9512 306892 9518
rect 306840 9454 306892 9460
rect 308036 9512 308088 9518
rect 308036 9454 308088 9460
rect 305920 9444 305972 9450
rect 305920 9386 305972 9392
rect 305828 8424 305880 8430
rect 305828 8366 305880 8372
rect 305552 4004 305604 4010
rect 305552 3946 305604 3952
rect 304908 3596 304960 3602
rect 304908 3538 304960 3544
rect 305564 480 305592 3946
rect 305932 3738 305960 9386
rect 306380 8424 306432 8430
rect 306380 8366 306432 8372
rect 305920 3732 305972 3738
rect 305920 3674 305972 3680
rect 306392 3534 306420 8366
rect 306748 4072 306800 4078
rect 306748 4014 306800 4020
rect 306380 3528 306432 3534
rect 306380 3470 306432 3476
rect 306760 480 306788 4014
rect 308048 3466 308076 9454
rect 308876 9314 308904 12022
rect 309888 9586 309916 12022
rect 309876 9580 309928 9586
rect 309876 9522 309928 9528
rect 308864 9308 308916 9314
rect 308864 9250 308916 9256
rect 310900 8838 310928 12022
rect 311820 9246 311848 12022
rect 311808 9240 311860 9246
rect 311808 9182 311860 9188
rect 312924 8906 312952 12022
rect 312912 8900 312964 8906
rect 312912 8842 312964 8848
rect 310888 8832 310940 8838
rect 310888 8774 310940 8780
rect 313936 8770 313964 12022
rect 314580 12022 314640 12050
rect 315652 12022 315896 12050
rect 316664 12022 317000 12050
rect 317676 12022 318012 12050
rect 314580 9178 314608 12022
rect 314568 9172 314620 9178
rect 314568 9114 314620 9120
rect 315868 9042 315896 12022
rect 316040 9580 316092 9586
rect 316040 9522 316092 9528
rect 316052 9382 316080 9522
rect 316040 9376 316092 9382
rect 316040 9318 316092 9324
rect 315856 9036 315908 9042
rect 315856 8978 315908 8984
rect 316972 8974 317000 12022
rect 317984 9450 318012 12022
rect 318628 12022 318688 12050
rect 319700 12022 320036 12050
rect 320712 12022 321048 12050
rect 321724 12022 322060 12050
rect 322736 12022 322888 12050
rect 323748 12022 324084 12050
rect 324760 12022 325096 12050
rect 325772 12022 326108 12050
rect 326784 12022 327028 12050
rect 327796 12022 328132 12050
rect 328808 12022 329144 12050
rect 317972 9444 318024 9450
rect 317972 9386 318024 9392
rect 316224 8968 316276 8974
rect 316224 8910 316276 8916
rect 316960 8968 317012 8974
rect 316960 8910 317012 8916
rect 313924 8764 313976 8770
rect 313924 8706 313976 8712
rect 310244 4140 310296 4146
rect 310244 4082 310296 4088
rect 309048 3868 309100 3874
rect 309048 3810 309100 3816
rect 307944 3460 307996 3466
rect 307944 3402 307996 3408
rect 308036 3460 308088 3466
rect 308036 3402 308088 3408
rect 307956 480 307984 3402
rect 309060 480 309088 3810
rect 310256 480 310284 4082
rect 311440 3936 311492 3942
rect 311440 3878 311492 3884
rect 311452 480 311480 3878
rect 312636 3800 312688 3806
rect 312636 3742 312688 3748
rect 312648 480 312676 3742
rect 313832 3664 313884 3670
rect 313832 3606 313884 3612
rect 313844 480 313872 3606
rect 315028 3596 315080 3602
rect 315028 3538 315080 3544
rect 315040 480 315068 3538
rect 316236 480 316264 8910
rect 318628 8702 318656 12022
rect 320008 9586 320036 12022
rect 319996 9580 320048 9586
rect 319996 9522 320048 9528
rect 321020 9518 321048 12022
rect 320916 9512 320968 9518
rect 320916 9454 320968 9460
rect 321008 9512 321060 9518
rect 321008 9454 321060 9460
rect 318616 8696 318668 8702
rect 318616 8638 318668 8644
rect 317328 3732 317380 3738
rect 317328 3674 317380 3680
rect 317340 480 317368 3674
rect 318524 3528 318576 3534
rect 318524 3470 318576 3476
rect 318536 480 318564 3470
rect 319720 3460 319772 3466
rect 319720 3402 319772 3408
rect 319732 480 319760 3402
rect 320928 480 320956 9454
rect 322032 9314 322060 12022
rect 322860 9654 322888 12022
rect 322848 9648 322900 9654
rect 322848 9590 322900 9596
rect 323308 9376 323360 9382
rect 323308 9318 323360 9324
rect 323400 9376 323452 9382
rect 323400 9318 323452 9324
rect 322020 9308 322072 9314
rect 322020 9250 322072 9256
rect 322112 9240 322164 9246
rect 322112 9182 322164 9188
rect 322124 480 322152 9182
rect 323320 480 323348 9318
rect 323412 8974 323440 9318
rect 323400 8968 323452 8974
rect 323400 8910 323452 8916
rect 323492 8968 323544 8974
rect 323492 8910 323544 8916
rect 323504 8702 323532 8910
rect 323492 8696 323544 8702
rect 323492 8638 323544 8644
rect 324056 8634 324084 12022
rect 325068 8838 325096 12022
rect 326080 9586 326108 12022
rect 326068 9580 326120 9586
rect 326068 9522 326120 9528
rect 325884 9512 325936 9518
rect 325884 9454 325936 9460
rect 325608 9172 325660 9178
rect 325608 9114 325660 9120
rect 324412 8832 324464 8838
rect 324412 8774 324464 8780
rect 325056 8832 325108 8838
rect 325056 8774 325108 8780
rect 324044 8628 324096 8634
rect 324044 8570 324096 8576
rect 324424 480 324452 8774
rect 325620 480 325648 9114
rect 325896 8498 325924 9454
rect 326804 8900 326856 8906
rect 326804 8842 326856 8848
rect 325884 8492 325936 8498
rect 325884 8434 325936 8440
rect 326816 480 326844 8842
rect 327000 8702 327028 12022
rect 328104 9518 328132 12022
rect 328000 9512 328052 9518
rect 328000 9454 328052 9460
rect 328092 9512 328144 9518
rect 328092 9454 328144 9460
rect 328012 9110 328040 9454
rect 327080 9104 327132 9110
rect 327080 9046 327132 9052
rect 328000 9104 328052 9110
rect 328000 9046 328052 9052
rect 326988 8696 327040 8702
rect 326988 8638 327040 8644
rect 327092 3126 327120 9046
rect 328000 8764 328052 8770
rect 328000 8706 328052 8712
rect 327080 3120 327132 3126
rect 327080 3062 327132 3068
rect 328012 480 328040 8706
rect 329116 8566 329144 12022
rect 329760 12022 329820 12050
rect 330832 12022 331168 12050
rect 331844 12022 332180 12050
rect 332856 12022 333192 12050
rect 329760 9246 329788 12022
rect 331036 9376 331088 9382
rect 331036 9318 331088 9324
rect 329748 9240 329800 9246
rect 329748 9182 329800 9188
rect 329656 9036 329708 9042
rect 329656 8978 329708 8984
rect 329104 8560 329156 8566
rect 329104 8502 329156 8508
rect 329668 3534 329696 8978
rect 330300 8628 330352 8634
rect 330300 8570 330352 8576
rect 329656 3528 329708 3534
rect 329656 3470 329708 3476
rect 330312 3398 330340 8570
rect 331048 6914 331076 9318
rect 331140 9178 331168 12022
rect 332152 9382 332180 12022
rect 332508 9444 332560 9450
rect 332508 9386 332560 9392
rect 332140 9376 332192 9382
rect 332140 9318 332192 9324
rect 331128 9172 331180 9178
rect 331128 9114 331180 9120
rect 331220 8968 331272 8974
rect 331220 8910 331272 8916
rect 331048 6886 331168 6914
rect 330392 3528 330444 3534
rect 330392 3470 330444 3476
rect 330300 3392 330352 3398
rect 330300 3334 330352 3340
rect 329196 3120 329248 3126
rect 329196 3062 329248 3068
rect 329208 480 329236 3062
rect 330404 480 330432 3470
rect 331140 2802 331168 6886
rect 331232 3602 331260 8910
rect 331220 3596 331272 3602
rect 331220 3538 331272 3544
rect 332520 3346 332548 9386
rect 332692 9104 332744 9110
rect 332692 9046 332744 9052
rect 332704 3466 332732 9046
rect 333164 8634 333192 12022
rect 333808 12022 333868 12050
rect 334880 12022 335216 12050
rect 335892 12022 336228 12050
rect 336904 12022 337240 12050
rect 337916 12022 338068 12050
rect 338928 12022 339264 12050
rect 339940 12022 340276 12050
rect 340952 12022 341288 12050
rect 341964 12022 342208 12050
rect 342976 12022 343312 12050
rect 343988 12022 344324 12050
rect 333808 9450 333836 12022
rect 334072 9512 334124 9518
rect 334072 9454 334124 9460
rect 333796 9444 333848 9450
rect 333796 9386 333848 9392
rect 333244 8832 333296 8838
rect 333244 8774 333296 8780
rect 333152 8628 333204 8634
rect 333152 8570 333204 8576
rect 333256 3534 333284 8774
rect 334084 3602 334112 9454
rect 335188 8838 335216 12022
rect 335544 9648 335596 9654
rect 335544 9590 335596 9596
rect 335452 9308 335504 9314
rect 335452 9250 335504 9256
rect 335176 8832 335228 8838
rect 335176 8774 335228 8780
rect 334164 8492 334216 8498
rect 334164 8434 334216 8440
rect 333888 3596 333940 3602
rect 333888 3538 333940 3544
rect 334072 3596 334124 3602
rect 334072 3538 334124 3544
rect 333244 3528 333296 3534
rect 333244 3470 333296 3476
rect 332692 3460 332744 3466
rect 332692 3402 332744 3408
rect 332520 3318 332732 3346
rect 331140 2774 331260 2802
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 354 331260 2774
rect 332704 480 332732 3318
rect 333900 480 333928 3538
rect 334176 3194 334204 8434
rect 335084 3460 335136 3466
rect 335084 3402 335136 3408
rect 334164 3188 334216 3194
rect 334164 3130 334216 3136
rect 335096 480 335124 3402
rect 335464 3126 335492 9250
rect 335556 3534 335584 9590
rect 336200 9110 336228 12022
rect 336188 9104 336240 9110
rect 336188 9046 336240 9052
rect 337212 8770 337240 12022
rect 338040 8906 338068 12022
rect 339236 8974 339264 12022
rect 340248 9654 340276 12022
rect 340236 9648 340288 9654
rect 340236 9590 340288 9596
rect 341260 9586 341288 12022
rect 340420 9580 340472 9586
rect 340420 9522 340472 9528
rect 341248 9580 341300 9586
rect 341248 9522 341300 9528
rect 339224 8968 339276 8974
rect 339224 8910 339276 8916
rect 338028 8900 338080 8906
rect 338028 8842 338080 8848
rect 337200 8764 337252 8770
rect 337200 8706 337252 8712
rect 335544 3528 335596 3534
rect 335544 3470 335596 3476
rect 338672 3528 338724 3534
rect 338672 3470 338724 3476
rect 336280 3188 336332 3194
rect 336280 3130 336332 3136
rect 335452 3120 335504 3126
rect 335452 3062 335504 3068
rect 336292 480 336320 3130
rect 337476 3120 337528 3126
rect 337476 3062 337528 3068
rect 337488 480 337516 3062
rect 338684 480 338712 3470
rect 339868 3392 339920 3398
rect 339868 3334 339920 3340
rect 339880 480 339908 3334
rect 340432 3058 340460 9522
rect 342180 8702 342208 12022
rect 343284 9518 343312 12022
rect 344296 9518 344324 12022
rect 344664 12022 345000 12050
rect 346012 12022 346348 12050
rect 347024 12022 347360 12050
rect 348036 12022 348372 12050
rect 343272 9512 343324 9518
rect 343272 9454 343324 9460
rect 343732 9512 343784 9518
rect 343732 9454 343784 9460
rect 344284 9512 344336 9518
rect 344284 9454 344336 9460
rect 343640 9308 343692 9314
rect 343640 9250 343692 9256
rect 340788 8696 340840 8702
rect 340788 8638 340840 8644
rect 342168 8696 342220 8702
rect 342168 8638 342220 8644
rect 340800 3194 340828 8638
rect 341984 8560 342036 8566
rect 341984 8502 342036 8508
rect 341996 3874 342024 8502
rect 341984 3868 342036 3874
rect 341984 3810 342036 3816
rect 343652 3466 343680 9250
rect 343744 3534 343772 9454
rect 344664 9314 344692 12022
rect 344652 9308 344704 9314
rect 344652 9250 344704 9256
rect 345204 9240 345256 9246
rect 345204 9182 345256 9188
rect 345216 3670 345244 9182
rect 346320 9042 346348 12022
rect 346584 9376 346636 9382
rect 346584 9318 346636 9324
rect 346492 9172 346544 9178
rect 346492 9114 346544 9120
rect 346308 9036 346360 9042
rect 346308 8978 346360 8984
rect 346400 8628 346452 8634
rect 346400 8570 346452 8576
rect 345756 3868 345808 3874
rect 345756 3810 345808 3816
rect 345204 3664 345256 3670
rect 345204 3606 345256 3612
rect 344560 3596 344612 3602
rect 344560 3538 344612 3544
rect 343732 3528 343784 3534
rect 343732 3470 343784 3476
rect 340972 3460 341024 3466
rect 340972 3402 341024 3408
rect 343640 3460 343692 3466
rect 343640 3402 343692 3408
rect 340788 3188 340840 3194
rect 340788 3130 340840 3136
rect 340420 3052 340472 3058
rect 340420 2994 340472 3000
rect 340984 480 341012 3402
rect 343364 3188 343416 3194
rect 343364 3130 343416 3136
rect 342168 3052 342220 3058
rect 342168 2994 342220 3000
rect 342180 480 342208 2994
rect 343376 480 343404 3130
rect 344572 480 344600 3538
rect 345768 480 345796 3810
rect 346412 3330 346440 8570
rect 346504 3602 346532 9114
rect 346492 3596 346544 3602
rect 346492 3538 346544 3544
rect 346596 3398 346624 9318
rect 347332 9314 347360 12022
rect 348344 9382 348372 12022
rect 348988 12022 349048 12050
rect 350060 12022 350396 12050
rect 351072 12022 351408 12050
rect 348332 9376 348384 9382
rect 348332 9318 348384 9324
rect 347320 9308 347372 9314
rect 347320 9250 347372 9256
rect 348988 8634 349016 12022
rect 350368 9450 350396 12022
rect 349068 9444 349120 9450
rect 349068 9386 349120 9392
rect 350356 9444 350408 9450
rect 350356 9386 350408 9392
rect 348976 8628 349028 8634
rect 348976 8570 349028 8576
rect 346952 3664 347004 3670
rect 346952 3606 347004 3612
rect 346584 3392 346636 3398
rect 346584 3334 346636 3340
rect 346400 3324 346452 3330
rect 346400 3266 346452 3272
rect 346964 480 346992 3606
rect 349080 3602 349108 9386
rect 351380 9246 351408 12022
rect 351932 12022 352084 12050
rect 352208 12022 353096 12050
rect 354108 12022 354444 12050
rect 355120 12022 355456 12050
rect 351368 9240 351420 9246
rect 351368 9182 351420 9188
rect 350540 8832 350592 8838
rect 350540 8774 350592 8780
rect 348056 3596 348108 3602
rect 348056 3538 348108 3544
rect 349068 3596 349120 3602
rect 349068 3538 349120 3544
rect 348068 480 348096 3538
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 349264 480 349292 3334
rect 350448 3324 350500 3330
rect 350448 3266 350500 3272
rect 350460 480 350488 3266
rect 350552 3058 350580 8774
rect 351932 3874 351960 12022
rect 352208 6914 352236 12022
rect 354416 9110 354444 12022
rect 354036 9104 354088 9110
rect 354036 9046 354088 9052
rect 354404 9104 354456 9110
rect 354404 9046 354456 9052
rect 353392 8900 353444 8906
rect 353392 8842 353444 8848
rect 353300 8764 353352 8770
rect 353300 8706 353352 8712
rect 352024 6886 352236 6914
rect 352024 6186 352052 6886
rect 352012 6180 352064 6186
rect 352012 6122 352064 6128
rect 351920 3868 351972 3874
rect 351920 3810 351972 3816
rect 353312 3602 353340 8706
rect 351644 3596 351696 3602
rect 351644 3538 351696 3544
rect 353300 3596 353352 3602
rect 353300 3538 353352 3544
rect 350540 3052 350592 3058
rect 350540 2994 350592 3000
rect 351656 480 351684 3538
rect 353404 3194 353432 8842
rect 353392 3188 353444 3194
rect 353392 3130 353444 3136
rect 352840 3052 352892 3058
rect 352840 2994 352892 3000
rect 352852 480 352880 2994
rect 354048 480 354076 9046
rect 355428 8906 355456 12022
rect 356072 12022 356132 12050
rect 356256 12022 357144 12050
rect 357452 12022 358156 12050
rect 359108 12022 359168 12050
rect 359292 12022 360180 12050
rect 361192 12022 361528 12050
rect 356072 9178 356100 12022
rect 356256 9466 356284 12022
rect 356336 9648 356388 9654
rect 356336 9590 356388 9596
rect 356164 9438 356284 9466
rect 356060 9172 356112 9178
rect 356060 9114 356112 9120
rect 356060 8968 356112 8974
rect 356060 8910 356112 8916
rect 355416 8900 355468 8906
rect 355416 8842 355468 8848
rect 355232 3596 355284 3602
rect 355232 3538 355284 3544
rect 355244 480 355272 3538
rect 356072 3534 356100 8910
rect 356164 3942 356192 9438
rect 356348 6914 356376 9590
rect 356256 6886 356376 6914
rect 356152 3936 356204 3942
rect 356152 3878 356204 3884
rect 356060 3528 356112 3534
rect 356060 3470 356112 3476
rect 356256 3058 356284 6886
rect 357452 3806 357480 12022
rect 358636 8696 358688 8702
rect 358636 8638 358688 8644
rect 357440 3800 357492 3806
rect 357440 3742 357492 3748
rect 357532 3528 357584 3534
rect 357532 3470 357584 3476
rect 356336 3188 356388 3194
rect 356336 3130 356388 3136
rect 356244 3052 356296 3058
rect 356244 2994 356296 3000
rect 356348 480 356376 3130
rect 357544 480 357572 3470
rect 358648 3126 358676 8638
rect 359108 8430 359136 12022
rect 359096 8424 359148 8430
rect 359096 8366 359148 8372
rect 359292 6914 359320 12022
rect 359924 9580 359976 9586
rect 359924 9522 359976 9528
rect 358924 6886 359320 6914
rect 358924 3738 358952 6886
rect 358912 3732 358964 3738
rect 358912 3674 358964 3680
rect 358636 3120 358688 3126
rect 358636 3062 358688 3068
rect 358728 3052 358780 3058
rect 358728 2994 358780 3000
rect 358740 480 358768 2994
rect 359936 480 359964 9522
rect 361500 8974 361528 12022
rect 361592 12022 362204 12050
rect 362972 12022 363216 12050
rect 363616 12022 364228 12050
rect 365240 12022 365576 12050
rect 366252 12022 366588 12050
rect 361488 8968 361540 8974
rect 361488 8910 361540 8916
rect 361592 6254 361620 12022
rect 361764 9512 361816 9518
rect 361764 9454 361816 9460
rect 361580 6248 361632 6254
rect 361580 6190 361632 6196
rect 361776 3534 361804 9454
rect 362224 8628 362276 8634
rect 362224 8570 362276 8576
rect 362236 4010 362264 8570
rect 362972 4146 363000 12022
rect 363616 6914 363644 12022
rect 365548 9246 365576 12022
rect 366560 9518 366588 12022
rect 367204 12022 367264 12050
rect 367480 12022 368276 12050
rect 369288 12022 369624 12050
rect 366548 9512 366600 9518
rect 366548 9454 366600 9460
rect 367008 9308 367060 9314
rect 367008 9250 367060 9256
rect 365444 9240 365496 9246
rect 365444 9182 365496 9188
rect 365536 9240 365588 9246
rect 365536 9182 365588 9188
rect 365456 8838 365484 9182
rect 365812 9036 365864 9042
rect 365812 8978 365864 8984
rect 365444 8832 365496 8838
rect 365444 8774 365496 8780
rect 364340 8424 364392 8430
rect 364340 8366 364392 8372
rect 363064 6886 363644 6914
rect 362960 4140 363012 4146
rect 362960 4082 363012 4088
rect 362224 4004 362276 4010
rect 362224 3946 362276 3952
rect 363064 3670 363092 6886
rect 364352 4962 364380 8366
rect 364340 4956 364392 4962
rect 364340 4898 364392 4904
rect 363052 3664 363104 3670
rect 363052 3606 363104 3612
rect 362316 3596 362368 3602
rect 362316 3538 362368 3544
rect 361764 3528 361816 3534
rect 361764 3470 361816 3476
rect 361120 3120 361172 3126
rect 361120 3062 361172 3068
rect 361132 480 361160 3062
rect 362328 480 362356 3538
rect 363512 3528 363564 3534
rect 363512 3470 363564 3476
rect 363524 480 363552 3470
rect 364616 3460 364668 3466
rect 364616 3402 364668 3408
rect 364628 480 364656 3402
rect 365824 480 365852 8978
rect 367020 480 367048 9250
rect 367204 3534 367232 12022
rect 367480 6914 367508 12022
rect 368296 9444 368348 9450
rect 368296 9386 368348 9392
rect 368204 9376 368256 9382
rect 368204 9318 368256 9324
rect 367296 6886 367508 6914
rect 367296 4894 367324 6886
rect 367284 4888 367336 4894
rect 367284 4830 367336 4836
rect 367192 3528 367244 3534
rect 367192 3470 367244 3476
rect 368216 480 368244 9318
rect 368308 3466 368336 9386
rect 369596 9042 369624 12022
rect 369872 12022 370300 12050
rect 371312 12022 371464 12050
rect 369584 9036 369636 9042
rect 369584 8978 369636 8984
rect 368388 8900 368440 8906
rect 368388 8842 368440 8848
rect 368400 3602 368428 8842
rect 369872 4010 369900 12022
rect 371436 9246 371464 12022
rect 371528 12022 372324 12050
rect 372632 12022 373336 12050
rect 374196 12022 374348 12050
rect 375208 12022 375360 12050
rect 375484 12022 376372 12050
rect 377384 12022 377628 12050
rect 370136 9240 370188 9246
rect 370136 9182 370188 9188
rect 371424 9240 371476 9246
rect 371424 9182 371476 9188
rect 370148 7614 370176 9182
rect 371148 8832 371200 8838
rect 371148 8774 371200 8780
rect 370136 7608 370188 7614
rect 370136 7550 370188 7556
rect 369400 4004 369452 4010
rect 369400 3946 369452 3952
rect 369860 4004 369912 4010
rect 369860 3946 369912 3952
rect 368388 3596 368440 3602
rect 368388 3538 368440 3544
rect 368296 3460 368348 3466
rect 368296 3402 368348 3408
rect 369412 480 369440 3946
rect 370596 3460 370648 3466
rect 370596 3402 370648 3408
rect 370608 480 370636 3402
rect 371160 2802 371188 8774
rect 371528 6914 371556 12022
rect 371884 9512 371936 9518
rect 371884 9454 371936 9460
rect 371252 6886 371556 6914
rect 371252 5030 371280 6886
rect 371896 6322 371924 9454
rect 371884 6316 371936 6322
rect 371884 6258 371936 6264
rect 371240 5024 371292 5030
rect 371240 4966 371292 4972
rect 372632 3466 372660 12022
rect 374196 6458 374224 12022
rect 375208 7750 375236 12022
rect 375288 9104 375340 9110
rect 375288 9046 375340 9052
rect 375196 7744 375248 7750
rect 375196 7686 375248 7692
rect 374184 6452 374236 6458
rect 374184 6394 374236 6400
rect 374092 6180 374144 6186
rect 374092 6122 374144 6128
rect 372896 3868 372948 3874
rect 372896 3810 372948 3816
rect 372620 3460 372672 3466
rect 372620 3402 372672 3408
rect 371160 2774 371280 2802
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 2774
rect 372908 480 372936 3810
rect 374104 480 374132 6122
rect 375196 3596 375248 3602
rect 375196 3538 375248 3544
rect 375208 3398 375236 3538
rect 375196 3392 375248 3398
rect 375196 3334 375248 3340
rect 375300 480 375328 9046
rect 375484 6914 375512 12022
rect 377600 7818 377628 12022
rect 378244 12022 378396 12050
rect 379072 12022 379408 12050
rect 379532 12022 380420 12050
rect 381432 12022 381768 12050
rect 378140 9512 378192 9518
rect 378140 9454 378192 9460
rect 377680 9172 377732 9178
rect 377680 9114 377732 9120
rect 377588 7812 377640 7818
rect 377588 7754 377640 7760
rect 375392 6886 375512 6914
rect 375392 4010 375420 6886
rect 375380 4004 375432 4010
rect 375380 3946 375432 3952
rect 376484 3392 376536 3398
rect 376484 3334 376536 3340
rect 376496 480 376524 3334
rect 377692 480 377720 9114
rect 378152 3534 378180 9454
rect 378244 6390 378272 12022
rect 379072 9518 379100 12022
rect 379060 9512 379112 9518
rect 379060 9454 379112 9460
rect 378232 6384 378284 6390
rect 378232 6326 378284 6332
rect 379532 4826 379560 12022
rect 381740 9110 381768 12022
rect 382384 12022 382444 12050
rect 383456 12022 383608 12050
rect 381728 9104 381780 9110
rect 381728 9046 381780 9052
rect 381176 4956 381228 4962
rect 381176 4898 381228 4904
rect 379520 4820 379572 4826
rect 379520 4762 379572 4768
rect 378876 3936 378928 3942
rect 378876 3878 378928 3884
rect 378140 3528 378192 3534
rect 378140 3470 378192 3476
rect 378888 480 378916 3878
rect 379980 3800 380032 3806
rect 379980 3742 380032 3748
rect 379992 480 380020 3742
rect 381188 480 381216 4898
rect 382384 4010 382412 12022
rect 383580 9178 383608 12022
rect 383672 12022 384468 12050
rect 385052 12022 385480 12050
rect 386432 12022 386492 12050
rect 386616 12022 387504 12050
rect 387812 12022 388516 12050
rect 389528 12022 389864 12050
rect 383568 9172 383620 9178
rect 383568 9114 383620 9120
rect 383568 8968 383620 8974
rect 383568 8910 383620 8916
rect 382372 4004 382424 4010
rect 382372 3946 382424 3952
rect 382372 3732 382424 3738
rect 382372 3674 382424 3680
rect 382384 480 382412 3674
rect 383580 480 383608 8910
rect 383672 4962 383700 12022
rect 384764 6248 384816 6254
rect 384764 6190 384816 6196
rect 383660 4956 383712 4962
rect 383660 4898 383712 4904
rect 384776 480 384804 6190
rect 385052 3806 385080 12022
rect 386432 7682 386460 12022
rect 386420 7676 386472 7682
rect 386420 7618 386472 7624
rect 386616 6914 386644 12022
rect 386432 6886 386644 6914
rect 386432 6186 386460 6886
rect 386420 6180 386472 6186
rect 386420 6122 386472 6128
rect 385960 4140 386012 4146
rect 385960 4082 386012 4088
rect 385040 3800 385092 3806
rect 385040 3742 385092 3748
rect 385972 480 386000 4082
rect 387812 3942 387840 12022
rect 389836 9314 389864 12022
rect 390480 12022 390540 12050
rect 390940 12022 391552 12050
rect 392044 12022 392564 12050
rect 393576 12022 393728 12050
rect 389824 9308 389876 9314
rect 389824 9250 389876 9256
rect 389732 9036 389784 9042
rect 389732 8978 389784 8984
rect 388260 7608 388312 7614
rect 388260 7550 388312 7556
rect 387800 3936 387852 3942
rect 387800 3878 387852 3884
rect 387156 3664 387208 3670
rect 387156 3606 387208 3612
rect 387168 480 387196 3606
rect 388272 480 388300 7550
rect 389456 6316 389508 6322
rect 389456 6258 389508 6264
rect 389468 480 389496 6258
rect 389744 5574 389772 8978
rect 390480 8974 390508 12022
rect 390468 8968 390520 8974
rect 390468 8910 390520 8916
rect 390940 6914 390968 12022
rect 391388 9240 391440 9246
rect 391388 9182 391440 9188
rect 390572 6886 390968 6914
rect 389732 5568 389784 5574
rect 389732 5510 389784 5516
rect 390572 4146 390600 6886
rect 391400 4350 391428 9182
rect 392044 6322 392072 12022
rect 393700 7614 393728 12022
rect 393792 12022 394588 12050
rect 394712 12022 395600 12050
rect 396092 12022 396612 12050
rect 397472 12022 397624 12050
rect 398636 12022 398788 12050
rect 393688 7608 393740 7614
rect 393688 7550 393740 7556
rect 393792 6914 393820 12022
rect 393332 6886 393820 6914
rect 392032 6316 392084 6322
rect 392032 6258 392084 6264
rect 393044 5568 393096 5574
rect 393044 5510 393096 5516
rect 391848 4888 391900 4894
rect 391848 4830 391900 4836
rect 391388 4344 391440 4350
rect 391388 4286 391440 4292
rect 390560 4140 390612 4146
rect 390560 4082 390612 4088
rect 390652 3596 390704 3602
rect 390652 3538 390704 3544
rect 390664 480 390692 3538
rect 391860 480 391888 4830
rect 393056 480 393084 5510
rect 393332 3670 393360 6886
rect 394712 4894 394740 12022
rect 396092 6254 396120 12022
rect 396080 6248 396132 6254
rect 396080 6190 396132 6196
rect 396540 5024 396592 5030
rect 396540 4966 396592 4972
rect 394700 4888 394752 4894
rect 394700 4830 394752 4836
rect 395344 4344 395396 4350
rect 395344 4286 395396 4292
rect 394240 4072 394292 4078
rect 394240 4014 394292 4020
rect 393320 3664 393372 3670
rect 393320 3606 393372 3612
rect 394252 480 394280 4014
rect 395356 480 395384 4286
rect 396552 480 396580 4966
rect 397472 3738 397500 12022
rect 398760 8906 398788 12022
rect 398852 12022 399648 12050
rect 400232 12022 400660 12050
rect 401672 12022 402008 12050
rect 402684 12022 402836 12050
rect 398748 8900 398800 8906
rect 398748 8842 398800 8848
rect 397460 3732 397512 3738
rect 397460 3674 397512 3680
rect 398852 3602 398880 12022
rect 400036 9172 400088 9178
rect 400036 9114 400088 9120
rect 400048 6526 400076 9114
rect 400128 7744 400180 7750
rect 400128 7686 400180 7692
rect 400036 6520 400088 6526
rect 400036 6462 400088 6468
rect 398932 6452 398984 6458
rect 398932 6394 398984 6400
rect 398840 3596 398892 3602
rect 398840 3538 398892 3544
rect 397736 3460 397788 3466
rect 397736 3402 397788 3408
rect 397748 480 397776 3402
rect 398944 480 398972 6394
rect 400140 480 400168 7686
rect 400232 3466 400260 12022
rect 401600 9104 401652 9110
rect 401600 9046 401652 9052
rect 400864 8900 400916 8906
rect 400864 8842 400916 8848
rect 400876 7954 400904 8842
rect 400864 7948 400916 7954
rect 400864 7890 400916 7896
rect 401612 7750 401640 9046
rect 401980 9042 402008 12022
rect 402808 9246 402836 12022
rect 402992 12022 403696 12050
rect 404708 12022 405044 12050
rect 402796 9240 402848 9246
rect 402796 9182 402848 9188
rect 401968 9036 402020 9042
rect 401968 8978 402020 8984
rect 402520 7812 402572 7818
rect 402520 7754 402572 7760
rect 401600 7744 401652 7750
rect 401600 7686 401652 7692
rect 401324 3868 401376 3874
rect 401324 3810 401376 3816
rect 400220 3460 400272 3466
rect 400220 3402 400272 3408
rect 401336 480 401364 3810
rect 402532 480 402560 7754
rect 402992 4078 403020 12022
rect 405016 9518 405044 12022
rect 405660 12022 405720 12050
rect 405844 12022 406732 12050
rect 407224 12022 407744 12050
rect 408696 12022 408756 12050
rect 408880 12022 409768 12050
rect 410780 12022 411116 12050
rect 405004 9512 405056 9518
rect 405004 9454 405056 9460
rect 403072 9308 403124 9314
rect 403072 9250 403124 9256
rect 403084 5098 403112 9250
rect 405660 9110 405688 12022
rect 405648 9104 405700 9110
rect 405648 9046 405700 9052
rect 405844 6914 405872 12022
rect 406384 9512 406436 9518
rect 406384 9454 406436 9460
rect 405752 6886 405872 6914
rect 403624 6384 403676 6390
rect 403624 6326 403676 6332
rect 403072 5092 403124 5098
rect 403072 5034 403124 5040
rect 402980 4072 403032 4078
rect 402980 4014 403032 4020
rect 403636 480 403664 6326
rect 405752 3874 405780 6886
rect 406396 5030 406424 9454
rect 407120 7744 407172 7750
rect 407120 7686 407172 7692
rect 406384 5024 406436 5030
rect 406384 4966 406436 4972
rect 406016 4820 406068 4826
rect 406016 4762 406068 4768
rect 405740 3868 405792 3874
rect 405740 3810 405792 3816
rect 404820 3528 404872 3534
rect 404820 3470 404872 3476
rect 404832 480 404860 3470
rect 406028 480 406056 4762
rect 407132 3482 407160 7686
rect 407224 6458 407252 12022
rect 408696 9518 408724 12022
rect 408684 9512 408736 9518
rect 408684 9454 408736 9460
rect 408880 6914 408908 12022
rect 411088 7886 411116 12022
rect 411272 12022 411792 12050
rect 412744 12022 412804 12050
rect 413816 12022 413968 12050
rect 414828 12022 415164 12050
rect 411168 9512 411220 9518
rect 411168 9454 411220 9460
rect 411076 7880 411128 7886
rect 411076 7822 411128 7828
rect 408512 6886 408908 6914
rect 407212 6452 407264 6458
rect 407212 6394 407264 6400
rect 408408 4004 408460 4010
rect 408408 3946 408460 3952
rect 407132 3454 407252 3482
rect 407224 480 407252 3454
rect 408420 480 408448 3946
rect 408512 3534 408540 6886
rect 409604 6520 409656 6526
rect 409604 6462 409656 6468
rect 408500 3528 408552 3534
rect 408500 3470 408552 3476
rect 409616 480 409644 6462
rect 411180 4962 411208 9454
rect 411272 6390 411300 12022
rect 411260 6384 411312 6390
rect 411260 6326 411312 6332
rect 410800 4956 410852 4962
rect 410800 4898 410852 4904
rect 411168 4956 411220 4962
rect 411168 4898 411220 4904
rect 410812 480 410840 4898
rect 412744 4010 412772 12022
rect 413940 9518 413968 12022
rect 413928 9512 413980 9518
rect 413928 9454 413980 9460
rect 415136 9382 415164 12022
rect 415412 12022 415840 12050
rect 416852 12022 417188 12050
rect 417864 12022 418108 12050
rect 418876 12022 419212 12050
rect 415124 9376 415176 9382
rect 415124 9318 415176 9324
rect 413836 8968 413888 8974
rect 413836 8910 413888 8916
rect 413848 8090 413876 8910
rect 413836 8084 413888 8090
rect 413836 8026 413888 8032
rect 413100 7744 413152 7750
rect 413100 7686 413152 7692
rect 412732 4004 412784 4010
rect 412732 3946 412784 3952
rect 411904 3800 411956 3806
rect 411904 3742 411956 3748
rect 411916 480 411944 3742
rect 413112 480 413140 7686
rect 414296 6180 414348 6186
rect 414296 6122 414348 6128
rect 414308 480 414336 6122
rect 415412 3806 415440 12022
rect 417160 7818 417188 12022
rect 417884 8084 417936 8090
rect 417884 8026 417936 8032
rect 417148 7812 417200 7818
rect 417148 7754 417200 7760
rect 416688 5092 416740 5098
rect 416688 5034 416740 5040
rect 415492 3936 415544 3942
rect 415492 3878 415544 3884
rect 415400 3800 415452 3806
rect 415400 3742 415452 3748
rect 415504 480 415532 3878
rect 416700 480 416728 5034
rect 417896 480 417924 8026
rect 418080 7750 418108 12022
rect 419184 9178 419212 12022
rect 419644 12022 419888 12050
rect 420840 12022 420900 12050
rect 421024 12022 421912 12050
rect 422312 12022 422924 12050
rect 423936 12022 424272 12050
rect 419356 9512 419408 9518
rect 419356 9454 419408 9460
rect 419172 9172 419224 9178
rect 419172 9114 419224 9120
rect 418804 9036 418856 9042
rect 418804 8978 418856 8984
rect 418068 7744 418120 7750
rect 418068 7686 418120 7692
rect 418816 6526 418844 8978
rect 418804 6520 418856 6526
rect 418804 6462 418856 6468
rect 419368 5166 419396 9454
rect 419644 6322 419672 12022
rect 420840 9042 420868 12022
rect 420828 9036 420880 9042
rect 420828 8978 420880 8984
rect 419540 6316 419592 6322
rect 419540 6258 419592 6264
rect 419632 6316 419684 6322
rect 419632 6258 419684 6264
rect 419552 5574 419580 6258
rect 419540 5568 419592 5574
rect 419540 5510 419592 5516
rect 420184 5568 420236 5574
rect 420184 5510 420236 5516
rect 419356 5160 419408 5166
rect 419356 5102 419408 5108
rect 418988 4140 419040 4146
rect 418988 4082 419040 4088
rect 419000 480 419028 4082
rect 420196 480 420224 5510
rect 421024 3942 421052 12022
rect 421472 9104 421524 9110
rect 421472 9046 421524 9052
rect 421484 7614 421512 9046
rect 421380 7608 421432 7614
rect 421380 7550 421432 7556
rect 421472 7608 421524 7614
rect 421472 7550 421524 7556
rect 421012 3936 421064 3942
rect 421012 3878 421064 3884
rect 421392 480 421420 7550
rect 422312 4826 422340 12022
rect 424244 9314 424272 12022
rect 424888 12022 424948 12050
rect 425960 12022 426296 12050
rect 424232 9308 424284 9314
rect 424232 9250 424284 9256
rect 424888 9110 424916 12022
rect 424876 9104 424928 9110
rect 424876 9046 424928 9052
rect 426268 7682 426296 12022
rect 426544 12022 426972 12050
rect 427832 12022 427984 12050
rect 428108 12022 428996 12050
rect 429212 12022 430008 12050
rect 431020 12022 431356 12050
rect 432032 12022 432184 12050
rect 426256 7676 426308 7682
rect 426256 7618 426308 7624
rect 426544 6254 426572 12022
rect 427268 7948 427320 7954
rect 427268 7890 427320 7896
rect 426532 6248 426584 6254
rect 426532 6190 426584 6196
rect 424968 6180 425020 6186
rect 424968 6122 425020 6128
rect 423772 4888 423824 4894
rect 423772 4830 423824 4836
rect 422300 4820 422352 4826
rect 422300 4762 422352 4768
rect 422576 3664 422628 3670
rect 422576 3606 422628 3612
rect 422588 480 422616 3606
rect 423784 480 423812 4830
rect 424980 480 425008 6122
rect 426164 3732 426216 3738
rect 426164 3674 426216 3680
rect 426176 480 426204 3674
rect 427280 480 427308 7890
rect 427832 3738 427860 12022
rect 428108 6914 428136 12022
rect 427924 6886 428136 6914
rect 427924 6186 427952 6886
rect 427912 6180 427964 6186
rect 427912 6122 427964 6128
rect 427820 3732 427872 3738
rect 427820 3674 427872 3680
rect 428464 3596 428516 3602
rect 428464 3538 428516 3544
rect 428476 480 428504 3538
rect 429212 3330 429240 12022
rect 430672 9376 430724 9382
rect 430672 9318 430724 9324
rect 430684 6594 430712 9318
rect 431328 8974 431356 12022
rect 432052 9512 432104 9518
rect 432052 9454 432104 9460
rect 431960 9240 432012 9246
rect 431960 9182 432012 9188
rect 431316 8968 431368 8974
rect 431316 8910 431368 8916
rect 430672 6588 430724 6594
rect 430672 6530 430724 6536
rect 430856 6520 430908 6526
rect 430856 6462 430908 6468
rect 429660 3460 429712 3466
rect 429660 3402 429712 3408
rect 429200 3324 429252 3330
rect 429200 3266 429252 3272
rect 429672 480 429700 3402
rect 430868 480 430896 6462
rect 431972 3074 432000 9182
rect 432064 3194 432092 9454
rect 432156 5098 432184 12022
rect 432708 12022 433044 12050
rect 433352 12022 434056 12050
rect 435008 12022 435068 12050
rect 435192 12022 436080 12050
rect 436296 12022 437092 12050
rect 437492 12022 438104 12050
rect 438872 12022 439116 12050
rect 439240 12022 440128 12050
rect 440344 12022 441140 12050
rect 441632 12022 442152 12050
rect 443012 12022 443164 12050
rect 443288 12022 444176 12050
rect 445188 12022 445524 12050
rect 432708 9518 432736 12022
rect 432696 9512 432748 9518
rect 432696 9454 432748 9460
rect 432144 5092 432196 5098
rect 432144 5034 432196 5040
rect 433248 4072 433300 4078
rect 433248 4014 433300 4020
rect 432052 3188 432104 3194
rect 432052 3130 432104 3136
rect 431972 3046 432092 3074
rect 432064 480 432092 3046
rect 433260 480 433288 4014
rect 433352 3602 433380 12022
rect 435008 7546 435036 12022
rect 434996 7540 435048 7546
rect 434996 7482 435048 7488
rect 435192 6914 435220 12022
rect 435548 7608 435600 7614
rect 435548 7550 435600 7556
rect 434732 6886 435220 6914
rect 434444 5024 434496 5030
rect 434444 4966 434496 4972
rect 433340 3596 433392 3602
rect 433340 3538 433392 3544
rect 434456 480 434484 4966
rect 434732 3670 434760 6886
rect 434720 3664 434772 3670
rect 434720 3606 434772 3612
rect 435560 480 435588 7550
rect 436296 6914 436324 12022
rect 436112 6886 436324 6914
rect 436112 3466 436140 6886
rect 437492 5030 437520 12022
rect 437940 6452 437992 6458
rect 437940 6394 437992 6400
rect 437480 5024 437532 5030
rect 437480 4966 437532 4972
rect 436744 3868 436796 3874
rect 436744 3810 436796 3816
rect 436100 3460 436152 3466
rect 436100 3402 436152 3408
rect 436756 480 436784 3810
rect 437952 480 437980 6394
rect 438872 3262 438900 12022
rect 439240 6914 439268 12022
rect 438964 6886 439268 6914
rect 438964 3398 438992 6886
rect 440344 6526 440372 12022
rect 441528 7880 441580 7886
rect 441528 7822 441580 7828
rect 440332 6520 440384 6526
rect 440332 6462 440384 6468
rect 439136 4956 439188 4962
rect 439136 4898 439188 4904
rect 438952 3392 439004 3398
rect 438952 3334 439004 3340
rect 438860 3256 438912 3262
rect 438860 3198 438912 3204
rect 439148 480 439176 4898
rect 440332 3528 440384 3534
rect 440332 3470 440384 3476
rect 440344 480 440372 3470
rect 441540 480 441568 7822
rect 441632 3534 441660 12022
rect 442632 6384 442684 6390
rect 442632 6326 442684 6332
rect 441620 3528 441672 3534
rect 441620 3470 441672 3476
rect 442644 480 442672 6326
rect 443012 4146 443040 12022
rect 443288 6914 443316 12022
rect 445496 9246 445524 12022
rect 445772 12022 446200 12050
rect 445668 9308 445720 9314
rect 445668 9250 445720 9256
rect 445484 9240 445536 9246
rect 445484 9182 445536 9188
rect 445680 7954 445708 9250
rect 445668 7948 445720 7954
rect 445668 7890 445720 7896
rect 443104 6886 443316 6914
rect 443104 4962 443132 6886
rect 445024 5160 445076 5166
rect 445024 5102 445076 5108
rect 443092 4956 443144 4962
rect 443092 4898 443144 4904
rect 443000 4140 443052 4146
rect 443000 4082 443052 4088
rect 443828 4004 443880 4010
rect 443828 3946 443880 3952
rect 443840 480 443868 3946
rect 445036 480 445064 5102
rect 445772 4078 445800 12022
rect 447198 11778 447226 12036
rect 447888 12022 448224 12050
rect 448532 12022 449236 12050
rect 450248 12022 450584 12050
rect 447198 11750 447272 11778
rect 447140 9512 447192 9518
rect 447140 9454 447192 9460
rect 446220 6588 446272 6594
rect 446220 6530 446272 6536
rect 445760 4072 445812 4078
rect 445760 4014 445812 4020
rect 446232 480 446260 6530
rect 447152 4894 447180 9454
rect 447244 6458 447272 11750
rect 447888 9518 447916 12022
rect 447876 9512 447928 9518
rect 447876 9454 447928 9460
rect 447232 6452 447284 6458
rect 447232 6394 447284 6400
rect 447140 4888 447192 4894
rect 447140 4830 447192 4836
rect 448532 4010 448560 12022
rect 450556 7886 450584 12022
rect 451200 12022 451260 12050
rect 451660 12022 452272 12050
rect 452764 12022 453284 12050
rect 454296 12022 454448 12050
rect 451200 9178 451228 12022
rect 450912 9172 450964 9178
rect 450912 9114 450964 9120
rect 451188 9172 451240 9178
rect 451188 9114 451240 9120
rect 450544 7880 450596 7886
rect 450544 7822 450596 7828
rect 448612 7812 448664 7818
rect 448612 7754 448664 7760
rect 448520 4004 448572 4010
rect 448520 3946 448572 3952
rect 447416 3800 447468 3806
rect 447416 3742 447468 3748
rect 447428 480 447456 3742
rect 448624 480 448652 7754
rect 449808 7744 449860 7750
rect 449808 7686 449860 7692
rect 449820 480 449848 7686
rect 450924 480 450952 9114
rect 451660 6914 451688 12022
rect 451292 6886 451688 6914
rect 451292 3874 451320 6886
rect 452764 6390 452792 12022
rect 454420 9518 454448 12022
rect 454512 12022 455308 12050
rect 456320 12022 456656 12050
rect 457332 12022 457668 12050
rect 454408 9512 454460 9518
rect 454408 9454 454460 9460
rect 453304 9036 453356 9042
rect 453304 8978 453356 8984
rect 452752 6384 452804 6390
rect 452752 6326 452804 6332
rect 452108 6316 452160 6322
rect 452108 6258 452160 6264
rect 451280 3868 451332 3874
rect 451280 3810 451332 3816
rect 452120 480 452148 6258
rect 453316 480 453344 8978
rect 454512 6914 454540 12022
rect 456628 7750 456656 12022
rect 456892 7948 456944 7954
rect 456892 7890 456944 7896
rect 456616 7744 456668 7750
rect 456616 7686 456668 7692
rect 454052 6886 454540 6914
rect 454052 3806 454080 6886
rect 455696 4820 455748 4826
rect 455696 4762 455748 4768
rect 454500 3936 454552 3942
rect 454500 3878 454552 3884
rect 454040 3800 454092 3806
rect 454040 3742 454092 3748
rect 454512 480 454540 3878
rect 455708 480 455736 4762
rect 456904 480 456932 7890
rect 457640 7818 457668 12022
rect 458192 12022 458344 12050
rect 459356 12022 459508 12050
rect 458088 9104 458140 9110
rect 458088 9046 458140 9052
rect 457628 7812 457680 7818
rect 457628 7754 457680 7760
rect 458100 480 458128 9046
rect 458192 3369 458220 12022
rect 459480 9450 459508 12022
rect 459664 12022 460368 12050
rect 460952 12022 461380 12050
rect 462392 12022 462728 12050
rect 463404 12022 463648 12050
rect 459468 9444 459520 9450
rect 459468 9386 459520 9392
rect 459192 7676 459244 7682
rect 459192 7618 459244 7624
rect 458178 3360 458234 3369
rect 458178 3295 458234 3304
rect 459204 480 459232 7618
rect 459664 6322 459692 12022
rect 459652 6316 459704 6322
rect 459652 6258 459704 6264
rect 460388 6248 460440 6254
rect 460388 6190 460440 6196
rect 460400 480 460428 6190
rect 460952 3942 460980 12022
rect 462700 8362 462728 12022
rect 463620 9382 463648 12022
rect 463712 12022 464416 12050
rect 465428 12022 465764 12050
rect 463608 9376 463660 9382
rect 463608 9318 463660 9324
rect 462688 8356 462740 8362
rect 462688 8298 462740 8304
rect 462780 6180 462832 6186
rect 462780 6122 462832 6128
rect 460940 3936 460992 3942
rect 460940 3878 460992 3884
rect 461584 3732 461636 3738
rect 461584 3674 461636 3680
rect 461596 480 461624 3674
rect 462792 480 462820 6122
rect 463712 3738 463740 12022
rect 465736 9314 465764 12022
rect 466380 12022 466440 12050
rect 467452 12022 467788 12050
rect 465724 9308 465776 9314
rect 465724 9250 465776 9256
rect 464068 9240 464120 9246
rect 464068 9182 464120 9188
rect 464080 5234 464108 9182
rect 466380 9110 466408 12022
rect 467196 9512 467248 9518
rect 467196 9454 467248 9460
rect 466368 9104 466420 9110
rect 466368 9046 466420 9052
rect 465172 8968 465224 8974
rect 465172 8910 465224 8916
rect 464068 5228 464120 5234
rect 464068 5170 464120 5176
rect 463700 3732 463752 3738
rect 463700 3674 463752 3680
rect 463976 3324 464028 3330
rect 463976 3266 464028 3272
rect 463988 480 464016 3266
rect 465184 480 465212 8910
rect 467208 5166 467236 9454
rect 467760 9042 467788 12022
rect 467852 12022 468464 12050
rect 469416 12022 469476 12050
rect 469600 12022 470488 12050
rect 471500 12022 471836 12050
rect 467748 9036 467800 9042
rect 467748 8978 467800 8984
rect 467852 6254 467880 12022
rect 469416 8566 469444 12022
rect 469404 8560 469456 8566
rect 469404 8502 469456 8508
rect 469600 6914 469628 12022
rect 471336 8560 471388 8566
rect 471336 8502 471388 8508
rect 469864 7608 469916 7614
rect 469864 7550 469916 7556
rect 469232 6886 469628 6914
rect 467840 6248 467892 6254
rect 467840 6190 467892 6196
rect 467196 5160 467248 5166
rect 467196 5102 467248 5108
rect 466276 5092 466328 5098
rect 466276 5034 466328 5040
rect 466288 480 466316 5034
rect 469232 3602 469260 6886
rect 468668 3596 468720 3602
rect 468668 3538 468720 3544
rect 469220 3596 469272 3602
rect 469220 3538 469272 3544
rect 467472 3188 467524 3194
rect 467472 3130 467524 3136
rect 467484 480 467512 3130
rect 468680 480 468708 3538
rect 469876 480 469904 7550
rect 471348 4826 471376 8502
rect 471808 7682 471836 12022
rect 471992 12022 472512 12050
rect 473524 12022 473860 12050
rect 474536 12022 474688 12050
rect 475548 12022 475884 12050
rect 471796 7676 471848 7682
rect 471796 7618 471848 7624
rect 471992 6186 472020 12022
rect 473832 8974 473860 12022
rect 474660 9246 474688 12022
rect 475856 9518 475884 12022
rect 476132 12022 476560 12050
rect 477572 12022 477908 12050
rect 478584 12022 478828 12050
rect 475844 9512 475896 9518
rect 475844 9454 475896 9460
rect 476028 9444 476080 9450
rect 476028 9386 476080 9392
rect 474648 9240 474700 9246
rect 474648 9182 474700 9188
rect 474096 9172 474148 9178
rect 474096 9114 474148 9120
rect 473820 8968 473872 8974
rect 473820 8910 473872 8916
rect 471980 6180 472032 6186
rect 471980 6122 472032 6128
rect 474108 5030 474136 9114
rect 476040 6730 476068 9386
rect 476028 6724 476080 6730
rect 476028 6666 476080 6672
rect 473452 5024 473504 5030
rect 473452 4966 473504 4972
rect 474096 5024 474148 5030
rect 474096 4966 474148 4972
rect 471336 4820 471388 4826
rect 471336 4762 471388 4768
rect 471060 3664 471112 3670
rect 471060 3606 471112 3612
rect 471072 480 471100 3606
rect 472256 3460 472308 3466
rect 472256 3402 472308 3408
rect 472268 480 472296 3402
rect 473464 480 473492 4966
rect 476132 3670 476160 12022
rect 477880 9450 477908 12022
rect 477868 9444 477920 9450
rect 477868 9386 477920 9392
rect 478800 7614 478828 12022
rect 478984 12022 479596 12050
rect 480272 12022 480608 12050
rect 481560 12022 481620 12050
rect 481744 12022 482632 12050
rect 483644 12022 483980 12050
rect 478880 9376 478932 9382
rect 478880 9318 478932 9324
rect 478788 7608 478840 7614
rect 478788 7550 478840 7556
rect 476948 6520 477000 6526
rect 476948 6462 477000 6468
rect 476120 3664 476172 3670
rect 476120 3606 476172 3612
rect 475752 3392 475804 3398
rect 475752 3334 475804 3340
rect 474556 3256 474608 3262
rect 474556 3198 474608 3204
rect 474568 480 474596 3198
rect 475764 480 475792 3334
rect 476960 480 476988 6462
rect 478892 5438 478920 9318
rect 478880 5432 478932 5438
rect 478880 5374 478932 5380
rect 478144 3528 478196 3534
rect 478144 3470 478196 3476
rect 478156 480 478184 3470
rect 478984 3466 479012 12022
rect 480272 5302 480300 12022
rect 481560 9178 481588 12022
rect 481548 9172 481600 9178
rect 481548 9114 481600 9120
rect 481744 6914 481772 12022
rect 483952 8090 483980 12022
rect 484412 12022 484656 12050
rect 485608 12022 485668 12050
rect 485792 12022 486680 12050
rect 487692 12022 488028 12050
rect 484308 9308 484360 9314
rect 484308 9250 484360 9256
rect 483940 8084 483992 8090
rect 483940 8026 483992 8032
rect 481652 6886 481772 6914
rect 480260 5296 480312 5302
rect 480260 5238 480312 5244
rect 480536 4956 480588 4962
rect 480536 4898 480588 4904
rect 479340 4140 479392 4146
rect 479340 4082 479392 4088
rect 478972 3460 479024 3466
rect 478972 3402 479024 3408
rect 479352 480 479380 4082
rect 480548 480 480576 4898
rect 481652 3534 481680 6886
rect 484320 6458 484348 9250
rect 484032 6452 484084 6458
rect 484032 6394 484084 6400
rect 484308 6452 484360 6458
rect 484308 6394 484360 6400
rect 481732 5228 481784 5234
rect 481732 5170 481784 5176
rect 481640 3528 481692 3534
rect 481640 3470 481692 3476
rect 481744 480 481772 5170
rect 482836 4072 482888 4078
rect 482836 4014 482888 4020
rect 482848 480 482876 4014
rect 484044 480 484072 6394
rect 484412 5370 484440 12022
rect 485136 9444 485188 9450
rect 485136 9386 485188 9392
rect 485148 6662 485176 9386
rect 485608 9314 485636 12022
rect 485596 9308 485648 9314
rect 485596 9250 485648 9256
rect 485136 6656 485188 6662
rect 485136 6598 485188 6604
rect 484400 5364 484452 5370
rect 484400 5306 484452 5312
rect 485792 5098 485820 12022
rect 488000 9450 488028 12022
rect 488552 12022 488704 12050
rect 488828 12022 489716 12050
rect 490728 12022 491064 12050
rect 491740 12022 492076 12050
rect 487988 9444 488040 9450
rect 487988 9386 488040 9392
rect 487620 7880 487672 7886
rect 487620 7822 487672 7828
rect 485780 5092 485832 5098
rect 485780 5034 485832 5040
rect 485228 4888 485280 4894
rect 485228 4830 485280 4836
rect 485240 480 485268 4830
rect 486424 4004 486476 4010
rect 486424 3946 486476 3952
rect 486436 480 486464 3946
rect 487632 480 487660 7822
rect 488552 3194 488580 12022
rect 488828 6914 488856 12022
rect 491036 8022 491064 12022
rect 492048 9654 492076 12022
rect 492692 12022 492752 12050
rect 492876 12022 493764 12050
rect 494072 12022 494776 12050
rect 495788 12022 496124 12050
rect 492036 9648 492088 9654
rect 492036 9590 492088 9596
rect 492588 9240 492640 9246
rect 492588 9182 492640 9188
rect 492600 8226 492628 9182
rect 492588 8220 492640 8226
rect 492588 8162 492640 8168
rect 491024 8016 491076 8022
rect 491024 7958 491076 7964
rect 488644 6886 488856 6914
rect 488644 5234 488672 6886
rect 491116 6384 491168 6390
rect 491116 6326 491168 6332
rect 488632 5228 488684 5234
rect 488632 5170 488684 5176
rect 488816 5024 488868 5030
rect 488816 4966 488868 4972
rect 488540 3188 488592 3194
rect 488540 3130 488592 3136
rect 488828 480 488856 4966
rect 489920 3868 489972 3874
rect 489920 3810 489972 3816
rect 489932 480 489960 3810
rect 491128 480 491156 6326
rect 492692 5166 492720 12022
rect 492876 6914 492904 12022
rect 492784 6886 492904 6914
rect 492784 6526 492812 6886
rect 492772 6520 492824 6526
rect 492772 6462 492824 6468
rect 492312 5160 492364 5166
rect 492312 5102 492364 5108
rect 492680 5160 492732 5166
rect 492680 5102 492732 5108
rect 492324 480 492352 5102
rect 493508 3800 493560 3806
rect 493508 3742 493560 3748
rect 493520 480 493548 3742
rect 494072 3262 494100 12022
rect 496096 9382 496124 12022
rect 496740 12022 496800 12050
rect 497812 12022 498148 12050
rect 498824 12022 499160 12050
rect 496740 9586 496768 12022
rect 496728 9580 496780 9586
rect 496728 9522 496780 9528
rect 496084 9376 496136 9382
rect 496084 9318 496136 9324
rect 498016 9376 498068 9382
rect 498016 9318 498068 9324
rect 495440 9104 495492 9110
rect 495440 9046 495492 9052
rect 495452 7886 495480 9046
rect 495440 7880 495492 7886
rect 495440 7822 495492 7828
rect 495900 7812 495952 7818
rect 495900 7754 495952 7760
rect 494704 7744 494756 7750
rect 494704 7686 494756 7692
rect 494060 3256 494112 3262
rect 494060 3198 494112 3204
rect 494716 480 494744 7686
rect 495912 480 495940 7754
rect 498028 6594 498056 9318
rect 498120 9110 498148 12022
rect 498200 9648 498252 9654
rect 498200 9590 498252 9596
rect 498212 9382 498240 9590
rect 498200 9376 498252 9382
rect 498200 9318 498252 9324
rect 498292 9172 498344 9178
rect 498292 9114 498344 9120
rect 498108 9104 498160 9110
rect 498108 9046 498160 9052
rect 498304 6730 498332 9114
rect 499132 7954 499160 12022
rect 499684 12022 499836 12050
rect 500512 12022 500848 12050
rect 501064 12022 501860 12050
rect 502872 12022 503208 12050
rect 503884 12022 504220 12050
rect 504896 12022 505048 12050
rect 505908 12022 506244 12050
rect 499580 9648 499632 9654
rect 499580 9590 499632 9596
rect 499120 7948 499172 7954
rect 499120 7890 499172 7896
rect 498200 6724 498252 6730
rect 498200 6666 498252 6672
rect 498292 6724 498344 6730
rect 498292 6666 498344 6672
rect 498016 6588 498068 6594
rect 498016 6530 498068 6536
rect 497094 3360 497150 3369
rect 497094 3295 497150 3304
rect 497108 480 497136 3295
rect 498212 480 498240 6666
rect 499396 6316 499448 6322
rect 499396 6258 499448 6264
rect 499408 480 499436 6258
rect 499592 4146 499620 9590
rect 499684 5030 499712 12022
rect 500512 9654 500540 12022
rect 500500 9648 500552 9654
rect 500500 9590 500552 9596
rect 501064 6390 501092 12022
rect 503180 9246 503208 12022
rect 503168 9240 503220 9246
rect 503168 9182 503220 9188
rect 504192 9178 504220 12022
rect 504916 9512 504968 9518
rect 504916 9454 504968 9460
rect 504180 9172 504232 9178
rect 504180 9114 504232 9120
rect 501788 8152 501840 8158
rect 501788 8094 501840 8100
rect 501052 6384 501104 6390
rect 501052 6326 501104 6332
rect 499672 5024 499724 5030
rect 499672 4966 499724 4972
rect 499580 4140 499632 4146
rect 499580 4082 499632 4088
rect 500592 3936 500644 3942
rect 500592 3878 500644 3884
rect 500604 480 500632 3878
rect 501800 480 501828 8094
rect 504928 6914 504956 9454
rect 505020 7750 505048 12022
rect 506216 7818 506244 12022
rect 506584 12022 506920 12050
rect 506480 7880 506532 7886
rect 506480 7822 506532 7828
rect 506204 7812 506256 7818
rect 506204 7754 506256 7760
rect 505008 7744 505060 7750
rect 505008 7686 505060 7692
rect 504928 6886 505048 6914
rect 505020 5438 505048 6886
rect 505376 6452 505428 6458
rect 505376 6394 505428 6400
rect 502984 5432 503036 5438
rect 502984 5374 503036 5380
rect 505008 5432 505060 5438
rect 505008 5374 505060 5380
rect 502996 480 503024 5374
rect 504180 3732 504232 3738
rect 504180 3674 504232 3680
rect 504192 480 504220 3674
rect 505388 480 505416 6394
rect 506492 480 506520 7822
rect 506584 3330 506612 12022
rect 507918 11778 507946 12036
rect 508056 12022 508944 12050
rect 509252 12022 509956 12050
rect 510908 12022 510968 12050
rect 511092 12022 511980 12050
rect 512104 12022 512992 12050
rect 513392 12022 514004 12050
rect 515016 12022 515168 12050
rect 507918 11750 507992 11778
rect 507676 9036 507728 9042
rect 507676 8978 507728 8984
rect 506572 3324 506624 3330
rect 506572 3266 506624 3272
rect 507688 480 507716 8978
rect 507964 6458 507992 11750
rect 507952 6452 508004 6458
rect 507952 6394 508004 6400
rect 508056 6322 508084 12022
rect 508044 6316 508096 6322
rect 508044 6258 508096 6264
rect 508872 6248 508924 6254
rect 508872 6190 508924 6196
rect 508884 480 508912 6190
rect 509252 3398 509280 12022
rect 510908 7886 510936 12022
rect 510896 7880 510948 7886
rect 510896 7822 510948 7828
rect 511092 6914 511120 12022
rect 512104 6914 512132 12022
rect 512460 7676 512512 7682
rect 512460 7618 512512 7624
rect 510632 6886 511120 6914
rect 512012 6886 512132 6914
rect 510632 4894 510660 6886
rect 510620 4888 510672 4894
rect 510620 4830 510672 4836
rect 510068 4820 510120 4826
rect 510068 4762 510120 4768
rect 509240 3392 509292 3398
rect 509240 3334 509292 3340
rect 510080 480 510108 4762
rect 512012 4010 512040 6886
rect 512000 4004 512052 4010
rect 512000 3946 512052 3952
rect 511264 3596 511316 3602
rect 511264 3538 511316 3544
rect 511276 480 511304 3538
rect 512472 480 512500 7618
rect 513392 4962 513420 12022
rect 515140 9042 515168 12022
rect 515232 12022 516028 12050
rect 516152 12022 517040 12050
rect 518052 12022 518388 12050
rect 515128 9036 515180 9042
rect 515128 8978 515180 8984
rect 514760 8968 514812 8974
rect 514760 8910 514812 8916
rect 513564 6180 513616 6186
rect 513564 6122 513616 6128
rect 513380 4956 513432 4962
rect 513380 4898 513432 4904
rect 513576 480 513604 6122
rect 514772 480 514800 8910
rect 515232 6914 515260 12022
rect 515956 8220 516008 8226
rect 515956 8162 516008 8168
rect 514864 6886 515260 6914
rect 514864 3942 514892 6886
rect 514852 3936 514904 3942
rect 514852 3878 514904 3884
rect 515968 480 515996 8162
rect 516152 6254 516180 12022
rect 518360 7682 518388 12022
rect 518912 12022 519064 12050
rect 520076 12022 520228 12050
rect 518348 7676 518400 7682
rect 518348 7618 518400 7624
rect 516140 6248 516192 6254
rect 516140 6190 516192 6196
rect 517152 5432 517204 5438
rect 517152 5374 517204 5380
rect 517164 480 517192 5374
rect 518912 4078 518940 12022
rect 520200 9518 520228 12022
rect 520384 12022 521088 12050
rect 521672 12022 522100 12050
rect 523052 12022 523112 12050
rect 523236 12022 524124 12050
rect 524432 12022 525136 12050
rect 526088 12022 526148 12050
rect 526272 12022 527160 12050
rect 527376 12022 528172 12050
rect 528572 12022 529184 12050
rect 529952 12022 530196 12050
rect 530320 12022 531208 12050
rect 531424 12022 532220 12050
rect 520188 9512 520240 9518
rect 520188 9454 520240 9460
rect 519636 9444 519688 9450
rect 519636 9386 519688 9392
rect 519648 6662 519676 9386
rect 519544 6656 519596 6662
rect 519544 6598 519596 6604
rect 519636 6656 519688 6662
rect 519636 6598 519688 6604
rect 518900 4072 518952 4078
rect 518900 4014 518952 4020
rect 518348 3664 518400 3670
rect 518348 3606 518400 3612
rect 518360 480 518388 3606
rect 519556 480 519584 6598
rect 520384 6186 520412 12022
rect 520740 7608 520792 7614
rect 520740 7550 520792 7556
rect 520372 6180 520424 6186
rect 520372 6122 520424 6128
rect 520752 480 520780 7550
rect 521672 3806 521700 12022
rect 523052 7614 523080 12022
rect 523040 7608 523092 7614
rect 523040 7550 523092 7556
rect 523236 6914 523264 12022
rect 523144 6886 523264 6914
rect 523040 5296 523092 5302
rect 523040 5238 523092 5244
rect 521660 3800 521712 3806
rect 521660 3742 521712 3748
rect 521844 3460 521896 3466
rect 521844 3402 521896 3408
rect 521856 480 521884 3402
rect 523052 480 523080 5238
rect 523144 4826 523172 6886
rect 524236 6724 524288 6730
rect 524236 6666 524288 6672
rect 523132 4820 523184 4826
rect 523132 4762 523184 4768
rect 524248 480 524276 6666
rect 524432 3874 524460 12022
rect 525432 9580 525484 9586
rect 525432 9522 525484 9528
rect 525444 5302 525472 9522
rect 526088 8974 526116 12022
rect 526076 8968 526128 8974
rect 526076 8910 526128 8916
rect 526272 6914 526300 12022
rect 526628 8084 526680 8090
rect 526628 8026 526680 8032
rect 525812 6886 526300 6914
rect 525432 5296 525484 5302
rect 525432 5238 525484 5244
rect 524420 3868 524472 3874
rect 524420 3810 524472 3816
rect 525812 3534 525840 6886
rect 525432 3528 525484 3534
rect 525432 3470 525484 3476
rect 525800 3528 525852 3534
rect 525800 3470 525852 3476
rect 525444 480 525472 3470
rect 526640 480 526668 8026
rect 527376 6914 527404 12022
rect 527192 6886 527404 6914
rect 527192 3670 527220 6886
rect 527824 5364 527876 5370
rect 527824 5306 527876 5312
rect 527180 3664 527232 3670
rect 527180 3606 527232 3612
rect 527836 480 527864 5306
rect 528572 3466 528600 12022
rect 529020 9308 529072 9314
rect 529020 9250 529072 9256
rect 528560 3460 528612 3466
rect 528560 3402 528612 3408
rect 529032 480 529060 9250
rect 529952 3738 529980 12022
rect 530320 6914 530348 12022
rect 530044 6886 530348 6914
rect 529940 3732 529992 3738
rect 529940 3674 529992 3680
rect 530044 3369 530072 6886
rect 531320 6656 531372 6662
rect 531320 6598 531372 6604
rect 530124 5092 530176 5098
rect 530124 5034 530176 5040
rect 530030 3360 530086 3369
rect 530030 3295 530086 3304
rect 530136 480 530164 5034
rect 531332 480 531360 6598
rect 531424 3602 531452 12022
rect 533436 9512 533488 9518
rect 533436 9454 533488 9460
rect 533448 5098 533476 9454
rect 536104 9376 536156 9382
rect 536104 9318 536156 9324
rect 534908 8016 534960 8022
rect 534908 7958 534960 7964
rect 533712 5228 533764 5234
rect 533712 5170 533764 5176
rect 533436 5092 533488 5098
rect 533436 5034 533488 5040
rect 531412 3596 531464 3602
rect 531412 3538 531464 3544
rect 532516 3188 532568 3194
rect 532516 3130 532568 3136
rect 532528 480 532556 3130
rect 533724 480 533752 5170
rect 534920 480 534948 7958
rect 536116 480 536144 9318
rect 546500 9240 546552 9246
rect 546500 9182 546552 9188
rect 543188 9104 543240 9110
rect 543188 9046 543240 9052
rect 540796 6588 540848 6594
rect 540796 6530 540848 6536
rect 538404 6520 538456 6526
rect 538404 6462 538456 6468
rect 537208 5160 537260 5166
rect 537208 5102 537260 5108
rect 537220 480 537248 5102
rect 538416 480 538444 6462
rect 539600 3256 539652 3262
rect 539600 3198 539652 3204
rect 539612 480 539640 3198
rect 540808 480 540836 6530
rect 541992 5296 542044 5302
rect 541992 5238 542044 5244
rect 542004 480 542032 5238
rect 543200 480 543228 9046
rect 544384 7948 544436 7954
rect 544384 7890 544436 7896
rect 544396 480 544424 7890
rect 545488 5024 545540 5030
rect 545488 4966 545540 4972
rect 545500 480 545528 4966
rect 546512 4690 546540 9182
rect 550272 9172 550324 9178
rect 550272 9114 550324 9120
rect 547880 6384 547932 6390
rect 547880 6326 547932 6332
rect 546500 4684 546552 4690
rect 546500 4626 546552 4632
rect 546684 4140 546736 4146
rect 546684 4082 546736 4088
rect 546696 480 546724 4082
rect 547892 480 547920 6326
rect 549076 4684 549128 4690
rect 549076 4626 549128 4632
rect 549088 480 549116 4626
rect 550284 480 550312 9114
rect 552664 7812 552716 7818
rect 552664 7754 552716 7760
rect 551468 7744 551520 7750
rect 551468 7686 551520 7692
rect 551480 480 551508 7686
rect 552676 480 552704 7754
rect 555436 6866 555464 19343
rect 563244 9036 563296 9042
rect 563244 8978 563296 8984
rect 558552 7880 558604 7886
rect 558552 7822 558604 7828
rect 555424 6860 555476 6866
rect 555424 6802 555476 6808
rect 554964 6452 555016 6458
rect 554964 6394 555016 6400
rect 553768 3324 553820 3330
rect 553768 3266 553820 3272
rect 553780 480 553808 3266
rect 554976 480 555004 6394
rect 556160 6316 556212 6322
rect 556160 6258 556212 6264
rect 556172 480 556200 6258
rect 557356 3392 557408 3398
rect 557356 3334 557408 3340
rect 557368 480 557396 3334
rect 558564 480 558592 7822
rect 562048 4956 562100 4962
rect 562048 4898 562100 4904
rect 559748 4888 559800 4894
rect 559748 4830 559800 4836
rect 559760 480 559788 4830
rect 560852 4004 560904 4010
rect 560852 3946 560904 3952
rect 560864 480 560892 3946
rect 562060 480 562088 4898
rect 563256 480 563284 8978
rect 576308 8968 576360 8974
rect 576308 8910 576360 8916
rect 566832 7676 566884 7682
rect 566832 7618 566884 7624
rect 565636 6248 565688 6254
rect 565636 6190 565688 6196
rect 564440 3936 564492 3942
rect 564440 3878 564492 3884
rect 564452 480 564480 3878
rect 565648 480 565676 6190
rect 566844 480 566872 7618
rect 572720 7608 572772 7614
rect 572720 7550 572772 7556
rect 570328 6180 570380 6186
rect 570328 6122 570380 6128
rect 569132 5092 569184 5098
rect 569132 5034 569184 5040
rect 568028 4072 568080 4078
rect 568028 4014 568080 4020
rect 568040 480 568068 4014
rect 569144 480 569172 5034
rect 570340 480 570368 6122
rect 571524 3800 571576 3806
rect 571524 3742 571576 3748
rect 571536 480 571564 3742
rect 572732 480 572760 7550
rect 573916 4820 573968 4826
rect 573916 4762 573968 4768
rect 573928 480 573956 4762
rect 575112 3868 575164 3874
rect 575112 3810 575164 3816
rect 575124 480 575152 3810
rect 576320 480 576348 8910
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581000 3732 581052 3738
rect 581000 3674 581052 3680
rect 578608 3664 578660 3670
rect 578608 3606 578660 3612
rect 577412 3528 577464 3534
rect 577412 3470 577464 3476
rect 577424 480 577452 3470
rect 578620 480 578648 3606
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 581012 480 581040 3674
rect 583392 3596 583444 3602
rect 583392 3538 583444 3544
rect 582194 3360 582250 3369
rect 582194 3295 582250 3304
rect 582208 480 582236 3295
rect 583404 480 583432 3538
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 697312 3478 697368
rect 3514 684256 3570 684312
rect 3422 645088 3478 645144
rect 3606 671200 3662 671256
rect 3514 632032 3570 632088
rect 580170 697176 580226 697232
rect 3698 658144 3754 658200
rect 580170 683848 580226 683904
rect 555422 655832 555478 655888
rect 9402 654744 9458 654800
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 555514 643592 555570 643648
rect 9402 642776 9458 642832
rect 580170 670656 580226 670692
rect 580262 657328 580318 657384
rect 580170 644000 580226 644056
rect 555606 631352 555662 631408
rect 9402 630808 9458 630864
rect 3606 619112 3662 619168
rect 3422 593000 3478 593056
rect 555146 619112 555202 619168
rect 9402 618840 9458 618896
rect 9402 606872 9458 606928
rect 3698 606056 3754 606112
rect 3514 579944 3570 580000
rect 3422 553832 3478 553888
rect 9402 594904 9458 594960
rect 555422 594632 555478 594688
rect 9402 582936 9458 582992
rect 8666 570968 8722 571024
rect 3606 566888 3662 566944
rect 3514 540776 3570 540832
rect 3422 514800 3478 514856
rect 9402 559000 9458 559056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 555698 606872 555754 606928
rect 580170 604152 580226 604208
rect 555514 582392 555570 582448
rect 555422 557912 555478 557968
rect 8666 547032 8722 547088
rect 9402 535064 9458 535120
rect 3606 527856 3662 527912
rect 9034 523096 9090 523152
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 555606 570152 555662 570208
rect 579802 564304 579858 564360
rect 555514 545672 555570 545728
rect 580170 551112 580226 551168
rect 580170 537784 580226 537840
rect 555606 533432 555662 533488
rect 555422 521192 555478 521248
rect 9402 511128 9458 511184
rect 3698 501744 3754 501800
rect 3514 488688 3570 488744
rect 9402 499160 9458 499216
rect 9034 487192 9090 487248
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 555698 508952 555754 509008
rect 580170 497936 580226 497992
rect 555514 496712 555570 496768
rect 555422 484472 555478 484528
rect 3606 475632 3662 475688
rect 3422 462576 3478 462632
rect 8666 475224 8722 475280
rect 9402 463256 9458 463312
rect 9034 451288 9090 451344
rect 3514 449520 3570 449576
rect 3422 436600 3478 436656
rect 580170 484608 580226 484664
rect 555606 472232 555662 472288
rect 579986 471416 580042 471472
rect 555514 459992 555570 460048
rect 580170 458088 580226 458144
rect 555422 447752 555478 447808
rect 9402 439320 9458 439376
rect 9402 427352 9458 427408
rect 3514 423544 3570 423600
rect 3422 410488 3478 410544
rect 580170 444760 580226 444816
rect 555514 435512 555570 435568
rect 580170 431568 580226 431624
rect 555422 423272 555478 423328
rect 9034 415384 9090 415440
rect 9402 403416 9458 403472
rect 580170 418240 580226 418296
rect 555514 411032 555570 411088
rect 580170 404912 580226 404968
rect 555422 398792 555478 398848
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3422 384376 3478 384432
rect 9402 391448 9458 391504
rect 7562 379480 7618 379536
rect 3422 371340 3478 371376
rect 3422 371320 3424 371340
rect 3424 371320 3476 371340
rect 3476 371320 3478 371340
rect 2962 358400 3018 358456
rect 3422 345364 3478 345400
rect 3422 345344 3424 345364
rect 3424 345344 3476 345364
rect 3476 345344 3478 345364
rect 580170 391720 580226 391776
rect 555514 386552 555570 386608
rect 580170 378392 580226 378448
rect 555422 374312 555478 374368
rect 9034 367512 9090 367568
rect 580170 365064 580226 365120
rect 555514 362072 555570 362128
rect 8942 355544 8998 355600
rect 3422 332308 3478 332344
rect 3422 332288 3424 332308
rect 3424 332288 3476 332308
rect 3476 332288 3478 332308
rect 9402 343596 9458 343632
rect 9402 343576 9404 343596
rect 9404 343576 9456 343596
rect 9456 343576 9458 343596
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 555606 349832 555662 349888
rect 580170 338544 580226 338600
rect 555422 337592 555478 337648
rect 8942 331608 8998 331664
rect 555514 325352 555570 325408
rect 580170 325216 580226 325272
rect 7562 319640 7618 319696
rect 3422 319232 3478 319288
rect 555422 313112 555478 313168
rect 580170 312024 580226 312080
rect 7654 307672 7710 307728
rect 2778 306176 2834 306232
rect 555514 300872 555570 300928
rect 580170 298696 580226 298752
rect 9494 295704 9550 295760
rect 2962 293120 3018 293176
rect 555422 288632 555478 288688
rect 580170 285368 580226 285424
rect 8666 283736 8722 283792
rect 3514 280064 3570 280120
rect 555422 276392 555478 276448
rect 579802 272176 579858 272232
rect 8206 271768 8262 271824
rect 3054 267144 3110 267200
rect 555422 264152 555478 264208
rect 9402 259800 9458 259856
rect 580170 258848 580226 258904
rect 3422 254108 3478 254144
rect 3422 254088 3424 254108
rect 3424 254088 3476 254108
rect 3476 254088 3478 254108
rect 556066 251912 556122 251968
rect 8942 247832 8998 247888
rect 579802 245520 579858 245576
rect 3698 241032 3754 241088
rect 555422 239672 555478 239728
rect 9402 235900 9404 235920
rect 9404 235900 9456 235920
rect 9456 235900 9458 235920
rect 9402 235864 9458 235900
rect 580170 232328 580226 232384
rect 4066 227976 4122 228032
rect 555422 227432 555478 227488
rect 8850 223896 8906 223952
rect 580170 219000 580226 219056
rect 555422 215192 555478 215248
rect 3146 214920 3202 214976
rect 9218 211928 9274 211984
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 555422 202952 555478 203008
rect 3422 201884 3478 201920
rect 3422 201864 3424 201884
rect 3424 201864 3476 201884
rect 3476 201864 3478 201884
rect 8298 199960 8354 200016
rect 580170 192480 580226 192536
rect 555422 190712 555478 190768
rect 3422 188808 3478 188864
rect 9402 187992 9458 188048
rect 580170 179152 580226 179208
rect 555422 178472 555478 178528
rect 9402 176024 9458 176080
rect 3330 175888 3386 175944
rect 555882 166268 555884 166288
rect 555884 166268 555936 166288
rect 555936 166268 555938 166288
rect 555882 166232 555938 166268
rect 580170 165824 580226 165880
rect 9402 164056 9458 164112
rect 3422 162868 3424 162888
rect 3424 162868 3476 162888
rect 3476 162868 3478 162888
rect 3422 162832 3478 162868
rect 555422 153992 555478 154048
rect 579526 152632 579582 152688
rect 8206 152088 8262 152144
rect 3422 149776 3478 149832
rect 555422 141752 555478 141808
rect 8206 140120 8262 140176
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 3238 136720 3294 136776
rect 555422 129512 555478 129568
rect 8206 128152 8262 128208
rect 580170 125976 580226 126032
rect 3422 123664 3478 123720
rect 555422 117272 555478 117328
rect 8942 116184 8998 116240
rect 579802 112784 579858 112840
rect 3422 110608 3478 110664
rect 555698 105032 555754 105088
rect 9402 104216 9458 104272
rect 4066 97552 4122 97608
rect 580170 99456 580226 99512
rect 554778 92792 554834 92848
rect 9402 92248 9458 92304
rect 4066 84632 4122 84688
rect 580170 86128 580226 86184
rect 555422 80552 555478 80608
rect 8942 80280 8998 80336
rect 580170 72936 580226 72992
rect 3422 71612 3424 71632
rect 3424 71612 3476 71632
rect 3476 71612 3478 71632
rect 3422 71576 3478 71612
rect 8942 68312 8998 68368
rect 555422 68312 555478 68368
rect 580170 59608 580226 59664
rect 3146 58520 3202 58576
rect 9402 56344 9458 56400
rect 555422 56072 555478 56128
rect 580170 46280 580226 46336
rect 2778 45500 2780 45520
rect 2780 45500 2832 45520
rect 2832 45500 2834 45520
rect 2778 45464 2834 45500
rect 9402 44376 9458 44432
rect 555422 43832 555478 43888
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 3422 32408 3478 32464
rect 9402 32408 9458 32464
rect 555514 31592 555570 31648
rect 9402 20440 9458 20496
rect 3514 19352 3570 19408
rect 579986 19760 580042 19816
rect 555422 19352 555478 19408
rect 3146 6468 3148 6488
rect 3148 6468 3200 6488
rect 3200 6468 3202 6488
rect 3146 6432 3202 6468
rect 39578 3304 39634 3360
rect 66258 3304 66314 3360
rect 78586 3304 78642 3360
rect 99746 3304 99802 3360
rect 458178 3304 458234 3360
rect 497094 3304 497150 3360
rect 530030 3304 530086 3360
rect 580170 6568 580226 6624
rect 582194 3304 582250 3360
<< metal3 >>
rect -960 697370 480 697460
rect 3417 697370 3483 697373
rect -960 697368 3483 697370
rect -960 697312 3422 697368
rect 3478 697312 3483 697368
rect -960 697310 3483 697312
rect -960 697220 480 697310
rect 3417 697307 3483 697310
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3509 684314 3575 684317
rect -960 684312 3575 684314
rect -960 684256 3514 684312
rect 3570 684256 3575 684312
rect -960 684254 3575 684256
rect -960 684164 480 684254
rect 3509 684251 3575 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3601 671258 3667 671261
rect -960 671256 3667 671258
rect -960 671200 3606 671256
rect 3662 671200 3667 671256
rect -960 671198 3667 671200
rect -960 671108 480 671198
rect 3601 671195 3667 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3693 658202 3759 658205
rect -960 658200 3759 658202
rect -960 658144 3698 658200
rect 3754 658144 3759 658200
rect -960 658142 3759 658144
rect -960 658052 480 658142
rect 3693 658139 3759 658142
rect 580257 657386 580323 657389
rect 583520 657386 584960 657476
rect 580257 657384 584960 657386
rect 580257 657328 580262 657384
rect 580318 657328 584960 657384
rect 580257 657326 584960 657328
rect 580257 657323 580323 657326
rect 583520 657236 584960 657326
rect 555417 655890 555483 655893
rect 553380 655888 555483 655890
rect 553380 655832 555422 655888
rect 555478 655832 555483 655888
rect 553380 655830 555483 655832
rect 555417 655827 555483 655830
rect 9397 654802 9463 654805
rect 9397 654800 12052 654802
rect 9397 654744 9402 654800
rect 9458 654744 12052 654800
rect 9397 654742 12052 654744
rect 9397 654739 9463 654742
rect -960 645146 480 645236
rect 3417 645146 3483 645149
rect -960 645144 3483 645146
rect -960 645088 3422 645144
rect 3478 645088 3483 645144
rect -960 645086 3483 645088
rect -960 644996 480 645086
rect 3417 645083 3483 645086
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 555509 643650 555575 643653
rect 553380 643648 555575 643650
rect 553380 643592 555514 643648
rect 555570 643592 555575 643648
rect 553380 643590 555575 643592
rect 555509 643587 555575 643590
rect 9397 642834 9463 642837
rect 9397 642832 12052 642834
rect 9397 642776 9402 642832
rect 9458 642776 12052 642832
rect 9397 642774 12052 642776
rect 9397 642771 9463 642774
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 555601 631410 555667 631413
rect 553380 631408 555667 631410
rect 553380 631352 555606 631408
rect 555662 631352 555667 631408
rect 553380 631350 555667 631352
rect 555601 631347 555667 631350
rect 9397 630866 9463 630869
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 9397 630864 12052 630866
rect 9397 630808 9402 630864
rect 9458 630808 12052 630864
rect 9397 630806 12052 630808
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 9397 630803 9463 630806
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3601 619170 3667 619173
rect 555141 619170 555207 619173
rect -960 619168 3667 619170
rect -960 619112 3606 619168
rect 3662 619112 3667 619168
rect -960 619110 3667 619112
rect 553380 619168 555207 619170
rect 553380 619112 555146 619168
rect 555202 619112 555207 619168
rect 553380 619110 555207 619112
rect -960 619020 480 619110
rect 3601 619107 3667 619110
rect 555141 619107 555207 619110
rect 9397 618898 9463 618901
rect 9397 618896 12052 618898
rect 9397 618840 9402 618896
rect 9458 618840 12052 618896
rect 9397 618838 12052 618840
rect 9397 618835 9463 618838
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 9397 606930 9463 606933
rect 555693 606930 555759 606933
rect 9397 606928 12052 606930
rect 9397 606872 9402 606928
rect 9458 606872 12052 606928
rect 9397 606870 12052 606872
rect 553380 606928 555759 606930
rect 553380 606872 555698 606928
rect 555754 606872 555759 606928
rect 553380 606870 555759 606872
rect 9397 606867 9463 606870
rect 555693 606867 555759 606870
rect -960 606114 480 606204
rect 3693 606114 3759 606117
rect -960 606112 3759 606114
rect -960 606056 3698 606112
rect 3754 606056 3759 606112
rect -960 606054 3759 606056
rect -960 605964 480 606054
rect 3693 606051 3759 606054
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect 9397 594962 9463 594965
rect 9397 594960 12052 594962
rect 9397 594904 9402 594960
rect 9458 594904 12052 594960
rect 9397 594902 12052 594904
rect 9397 594899 9463 594902
rect 555417 594690 555483 594693
rect 553380 594688 555483 594690
rect 553380 594632 555422 594688
rect 555478 594632 555483 594688
rect 553380 594630 555483 594632
rect 555417 594627 555483 594630
rect -960 593058 480 593148
rect 3417 593058 3483 593061
rect -960 593056 3483 593058
rect -960 593000 3422 593056
rect 3478 593000 3483 593056
rect -960 592998 3483 593000
rect -960 592908 480 592998
rect 3417 592995 3483 592998
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 9397 582994 9463 582997
rect 9397 582992 12052 582994
rect 9397 582936 9402 582992
rect 9458 582936 12052 582992
rect 9397 582934 12052 582936
rect 9397 582931 9463 582934
rect 555509 582450 555575 582453
rect 553380 582448 555575 582450
rect 553380 582392 555514 582448
rect 555570 582392 555575 582448
rect 553380 582390 555575 582392
rect 555509 582387 555575 582390
rect -960 580002 480 580092
rect 3509 580002 3575 580005
rect -960 580000 3575 580002
rect -960 579944 3514 580000
rect 3570 579944 3575 580000
rect -960 579942 3575 579944
rect -960 579852 480 579942
rect 3509 579939 3575 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 8661 571026 8727 571029
rect 8661 571024 12052 571026
rect 8661 570968 8666 571024
rect 8722 570968 12052 571024
rect 8661 570966 12052 570968
rect 8661 570963 8727 570966
rect 555601 570210 555667 570213
rect 553380 570208 555667 570210
rect 553380 570152 555606 570208
rect 555662 570152 555667 570208
rect 553380 570150 555667 570152
rect 555601 570147 555667 570150
rect -960 566946 480 567036
rect 3601 566946 3667 566949
rect -960 566944 3667 566946
rect -960 566888 3606 566944
rect 3662 566888 3667 566944
rect -960 566886 3667 566888
rect -960 566796 480 566886
rect 3601 566883 3667 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect 9397 559058 9463 559061
rect 9397 559056 12052 559058
rect 9397 559000 9402 559056
rect 9458 559000 12052 559056
rect 9397 558998 12052 559000
rect 9397 558995 9463 558998
rect 555417 557970 555483 557973
rect 553380 557968 555483 557970
rect 553380 557912 555422 557968
rect 555478 557912 555483 557968
rect 553380 557910 555483 557912
rect 555417 557907 555483 557910
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 580165 551170 580231 551173
rect 583520 551170 584960 551260
rect 580165 551168 584960 551170
rect 580165 551112 580170 551168
rect 580226 551112 584960 551168
rect 580165 551110 584960 551112
rect 580165 551107 580231 551110
rect 583520 551020 584960 551110
rect 8661 547090 8727 547093
rect 8661 547088 12052 547090
rect 8661 547032 8666 547088
rect 8722 547032 12052 547088
rect 8661 547030 12052 547032
rect 8661 547027 8727 547030
rect 555509 545730 555575 545733
rect 553380 545728 555575 545730
rect 553380 545672 555514 545728
rect 555570 545672 555575 545728
rect 553380 545670 555575 545672
rect 555509 545667 555575 545670
rect -960 540834 480 540924
rect 3509 540834 3575 540837
rect -960 540832 3575 540834
rect -960 540776 3514 540832
rect 3570 540776 3575 540832
rect -960 540774 3575 540776
rect -960 540684 480 540774
rect 3509 540771 3575 540774
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 9397 535122 9463 535125
rect 9397 535120 12052 535122
rect 9397 535064 9402 535120
rect 9458 535064 12052 535120
rect 9397 535062 12052 535064
rect 9397 535059 9463 535062
rect 555601 533490 555667 533493
rect 553380 533488 555667 533490
rect 553380 533432 555606 533488
rect 555662 533432 555667 533488
rect 553380 533430 555667 533432
rect 555601 533427 555667 533430
rect -960 527914 480 528004
rect 3601 527914 3667 527917
rect -960 527912 3667 527914
rect -960 527856 3606 527912
rect 3662 527856 3667 527912
rect -960 527854 3667 527856
rect -960 527764 480 527854
rect 3601 527851 3667 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 9029 523154 9095 523157
rect 9029 523152 12052 523154
rect 9029 523096 9034 523152
rect 9090 523096 12052 523152
rect 9029 523094 12052 523096
rect 9029 523091 9095 523094
rect 555417 521250 555483 521253
rect 553380 521248 555483 521250
rect 553380 521192 555422 521248
rect 555478 521192 555483 521248
rect 553380 521190 555483 521192
rect 555417 521187 555483 521190
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 9397 511186 9463 511189
rect 9397 511184 12052 511186
rect 9397 511128 9402 511184
rect 9458 511128 12052 511184
rect 583520 511172 584960 511262
rect 9397 511126 12052 511128
rect 9397 511123 9463 511126
rect 555693 509010 555759 509013
rect 553380 509008 555759 509010
rect 553380 508952 555698 509008
rect 555754 508952 555759 509008
rect 553380 508950 555759 508952
rect 555693 508947 555759 508950
rect -960 501802 480 501892
rect 3693 501802 3759 501805
rect -960 501800 3759 501802
rect -960 501744 3698 501800
rect 3754 501744 3759 501800
rect -960 501742 3759 501744
rect -960 501652 480 501742
rect 3693 501739 3759 501742
rect 9397 499218 9463 499221
rect 9397 499216 12052 499218
rect 9397 499160 9402 499216
rect 9458 499160 12052 499216
rect 9397 499158 12052 499160
rect 9397 499155 9463 499158
rect 580165 497994 580231 497997
rect 583520 497994 584960 498084
rect 580165 497992 584960 497994
rect 580165 497936 580170 497992
rect 580226 497936 584960 497992
rect 580165 497934 584960 497936
rect 580165 497931 580231 497934
rect 583520 497844 584960 497934
rect 555509 496770 555575 496773
rect 553380 496768 555575 496770
rect 553380 496712 555514 496768
rect 555570 496712 555575 496768
rect 553380 496710 555575 496712
rect 555509 496707 555575 496710
rect -960 488746 480 488836
rect 3509 488746 3575 488749
rect -960 488744 3575 488746
rect -960 488688 3514 488744
rect 3570 488688 3575 488744
rect -960 488686 3575 488688
rect -960 488596 480 488686
rect 3509 488683 3575 488686
rect 9029 487250 9095 487253
rect 9029 487248 12052 487250
rect 9029 487192 9034 487248
rect 9090 487192 12052 487248
rect 9029 487190 12052 487192
rect 9029 487187 9095 487190
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 555417 484530 555483 484533
rect 553380 484528 555483 484530
rect 553380 484472 555422 484528
rect 555478 484472 555483 484528
rect 583520 484516 584960 484606
rect 553380 484470 555483 484472
rect 555417 484467 555483 484470
rect -960 475690 480 475780
rect 3601 475690 3667 475693
rect -960 475688 3667 475690
rect -960 475632 3606 475688
rect 3662 475632 3667 475688
rect -960 475630 3667 475632
rect -960 475540 480 475630
rect 3601 475627 3667 475630
rect 8661 475282 8727 475285
rect 8661 475280 12052 475282
rect 8661 475224 8666 475280
rect 8722 475224 12052 475280
rect 8661 475222 12052 475224
rect 8661 475219 8727 475222
rect 555601 472290 555667 472293
rect 553380 472288 555667 472290
rect 553380 472232 555606 472288
rect 555662 472232 555667 472288
rect 553380 472230 555667 472232
rect 555601 472227 555667 472230
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 9397 463314 9463 463317
rect 9397 463312 12052 463314
rect 9397 463256 9402 463312
rect 9458 463256 12052 463312
rect 9397 463254 12052 463256
rect 9397 463251 9463 463254
rect -960 462634 480 462724
rect 3417 462634 3483 462637
rect -960 462632 3483 462634
rect -960 462576 3422 462632
rect 3478 462576 3483 462632
rect -960 462574 3483 462576
rect -960 462484 480 462574
rect 3417 462571 3483 462574
rect 555509 460050 555575 460053
rect 553380 460048 555575 460050
rect 553380 459992 555514 460048
rect 555570 459992 555575 460048
rect 553380 459990 555575 459992
rect 555509 459987 555575 459990
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 9029 451346 9095 451349
rect 9029 451344 12052 451346
rect 9029 451288 9034 451344
rect 9090 451288 12052 451344
rect 9029 451286 12052 451288
rect 9029 451283 9095 451286
rect -960 449578 480 449668
rect 3509 449578 3575 449581
rect -960 449576 3575 449578
rect -960 449520 3514 449576
rect 3570 449520 3575 449576
rect -960 449518 3575 449520
rect -960 449428 480 449518
rect 3509 449515 3575 449518
rect 555417 447810 555483 447813
rect 553380 447808 555483 447810
rect 553380 447752 555422 447808
rect 555478 447752 555483 447808
rect 553380 447750 555483 447752
rect 555417 447747 555483 447750
rect 580165 444818 580231 444821
rect 583520 444818 584960 444908
rect 580165 444816 584960 444818
rect 580165 444760 580170 444816
rect 580226 444760 584960 444816
rect 580165 444758 584960 444760
rect 580165 444755 580231 444758
rect 583520 444668 584960 444758
rect 9397 439378 9463 439381
rect 9397 439376 12052 439378
rect 9397 439320 9402 439376
rect 9458 439320 12052 439376
rect 9397 439318 12052 439320
rect 9397 439315 9463 439318
rect -960 436658 480 436748
rect 3417 436658 3483 436661
rect -960 436656 3483 436658
rect -960 436600 3422 436656
rect 3478 436600 3483 436656
rect -960 436598 3483 436600
rect -960 436508 480 436598
rect 3417 436595 3483 436598
rect 555509 435570 555575 435573
rect 553380 435568 555575 435570
rect 553380 435512 555514 435568
rect 555570 435512 555575 435568
rect 553380 435510 555575 435512
rect 555509 435507 555575 435510
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 9397 427410 9463 427413
rect 9397 427408 12052 427410
rect 9397 427352 9402 427408
rect 9458 427352 12052 427408
rect 9397 427350 12052 427352
rect 9397 427347 9463 427350
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 555417 423330 555483 423333
rect 553380 423328 555483 423330
rect 553380 423272 555422 423328
rect 555478 423272 555483 423328
rect 553380 423270 555483 423272
rect 555417 423267 555483 423270
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 9029 415442 9095 415445
rect 9029 415440 12052 415442
rect 9029 415384 9034 415440
rect 9090 415384 12052 415440
rect 9029 415382 12052 415384
rect 9029 415379 9095 415382
rect 555509 411090 555575 411093
rect 553380 411088 555575 411090
rect 553380 411032 555514 411088
rect 555570 411032 555575 411088
rect 553380 411030 555575 411032
rect 555509 411027 555575 411030
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 9397 403474 9463 403477
rect 9397 403472 12052 403474
rect 9397 403416 9402 403472
rect 9458 403416 12052 403472
rect 9397 403414 12052 403416
rect 9397 403411 9463 403414
rect 555417 398850 555483 398853
rect 553380 398848 555483 398850
rect 553380 398792 555422 398848
rect 555478 398792 555483 398848
rect 553380 398790 555483 398792
rect 555417 398787 555483 398790
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 580165 391778 580231 391781
rect 583520 391778 584960 391868
rect 580165 391776 584960 391778
rect 580165 391720 580170 391776
rect 580226 391720 584960 391776
rect 580165 391718 584960 391720
rect 580165 391715 580231 391718
rect 583520 391628 584960 391718
rect 9397 391506 9463 391509
rect 9397 391504 12052 391506
rect 9397 391448 9402 391504
rect 9458 391448 12052 391504
rect 9397 391446 12052 391448
rect 9397 391443 9463 391446
rect 555509 386610 555575 386613
rect 553380 386608 555575 386610
rect 553380 386552 555514 386608
rect 555570 386552 555575 386608
rect 553380 386550 555575 386552
rect 555509 386547 555575 386550
rect -960 384434 480 384524
rect 3417 384434 3483 384437
rect -960 384432 3483 384434
rect -960 384376 3422 384432
rect 3478 384376 3483 384432
rect -960 384374 3483 384376
rect -960 384284 480 384374
rect 3417 384371 3483 384374
rect 7557 379538 7623 379541
rect 7557 379536 12052 379538
rect 7557 379480 7562 379536
rect 7618 379480 12052 379536
rect 7557 379478 12052 379480
rect 7557 379475 7623 379478
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 555417 374370 555483 374373
rect 553380 374368 555483 374370
rect 553380 374312 555422 374368
rect 555478 374312 555483 374368
rect 553380 374310 555483 374312
rect 555417 374307 555483 374310
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 9029 367570 9095 367573
rect 9029 367568 12052 367570
rect 9029 367512 9034 367568
rect 9090 367512 12052 367568
rect 9029 367510 12052 367512
rect 9029 367507 9095 367510
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 555509 362130 555575 362133
rect 553380 362128 555575 362130
rect 553380 362072 555514 362128
rect 555570 362072 555575 362128
rect 553380 362070 555575 362072
rect 555509 362067 555575 362070
rect -960 358458 480 358548
rect 2957 358458 3023 358461
rect -960 358456 3023 358458
rect -960 358400 2962 358456
rect 3018 358400 3023 358456
rect -960 358398 3023 358400
rect -960 358308 480 358398
rect 2957 358395 3023 358398
rect 8937 355602 9003 355605
rect 8937 355600 12052 355602
rect 8937 355544 8942 355600
rect 8998 355544 12052 355600
rect 8937 355542 12052 355544
rect 8937 355539 9003 355542
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 555601 349890 555667 349893
rect 553380 349888 555667 349890
rect 553380 349832 555606 349888
rect 555662 349832 555667 349888
rect 553380 349830 555667 349832
rect 555601 349827 555667 349830
rect -960 345402 480 345492
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 9397 343634 9463 343637
rect 9397 343632 12052 343634
rect 9397 343576 9402 343632
rect 9458 343576 12052 343632
rect 9397 343574 12052 343576
rect 9397 343571 9463 343574
rect 580165 338602 580231 338605
rect 583520 338602 584960 338692
rect 580165 338600 584960 338602
rect 580165 338544 580170 338600
rect 580226 338544 584960 338600
rect 580165 338542 584960 338544
rect 580165 338539 580231 338542
rect 583520 338452 584960 338542
rect 555417 337650 555483 337653
rect 553380 337648 555483 337650
rect 553380 337592 555422 337648
rect 555478 337592 555483 337648
rect 553380 337590 555483 337592
rect 555417 337587 555483 337590
rect -960 332346 480 332436
rect 3417 332346 3483 332349
rect -960 332344 3483 332346
rect -960 332288 3422 332344
rect 3478 332288 3483 332344
rect -960 332286 3483 332288
rect -960 332196 480 332286
rect 3417 332283 3483 332286
rect 8937 331666 9003 331669
rect 8937 331664 12052 331666
rect 8937 331608 8942 331664
rect 8998 331608 12052 331664
rect 8937 331606 12052 331608
rect 8937 331603 9003 331606
rect 555509 325410 555575 325413
rect 553380 325408 555575 325410
rect 553380 325352 555514 325408
rect 555570 325352 555575 325408
rect 553380 325350 555575 325352
rect 555509 325347 555575 325350
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 7557 319698 7623 319701
rect 7557 319696 12052 319698
rect 7557 319640 7562 319696
rect 7618 319640 12052 319696
rect 7557 319638 12052 319640
rect 7557 319635 7623 319638
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 555417 313170 555483 313173
rect 553380 313168 555483 313170
rect 553380 313112 555422 313168
rect 555478 313112 555483 313168
rect 553380 313110 555483 313112
rect 555417 313107 555483 313110
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 7649 307730 7715 307733
rect 7649 307728 12052 307730
rect 7649 307672 7654 307728
rect 7710 307672 12052 307728
rect 7649 307670 12052 307672
rect 7649 307667 7715 307670
rect -960 306234 480 306324
rect 2773 306234 2839 306237
rect -960 306232 2839 306234
rect -960 306176 2778 306232
rect 2834 306176 2839 306232
rect -960 306174 2839 306176
rect -960 306084 480 306174
rect 2773 306171 2839 306174
rect 555509 300930 555575 300933
rect 553380 300928 555575 300930
rect 553380 300872 555514 300928
rect 555570 300872 555575 300928
rect 553380 300870 555575 300872
rect 555509 300867 555575 300870
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 9489 295762 9555 295765
rect 9489 295760 12052 295762
rect 9489 295704 9494 295760
rect 9550 295704 12052 295760
rect 9489 295702 12052 295704
rect 9489 295699 9555 295702
rect -960 293178 480 293268
rect 2957 293178 3023 293181
rect -960 293176 3023 293178
rect -960 293120 2962 293176
rect 3018 293120 3023 293176
rect -960 293118 3023 293120
rect -960 293028 480 293118
rect 2957 293115 3023 293118
rect 555417 288690 555483 288693
rect 553380 288688 555483 288690
rect 553380 288632 555422 288688
rect 555478 288632 555483 288688
rect 553380 288630 555483 288632
rect 555417 288627 555483 288630
rect 580165 285426 580231 285429
rect 583520 285426 584960 285516
rect 580165 285424 584960 285426
rect 580165 285368 580170 285424
rect 580226 285368 584960 285424
rect 580165 285366 584960 285368
rect 580165 285363 580231 285366
rect 583520 285276 584960 285366
rect 8661 283794 8727 283797
rect 8661 283792 12052 283794
rect 8661 283736 8666 283792
rect 8722 283736 12052 283792
rect 8661 283734 12052 283736
rect 8661 283731 8727 283734
rect -960 280122 480 280212
rect 3509 280122 3575 280125
rect -960 280120 3575 280122
rect -960 280064 3514 280120
rect 3570 280064 3575 280120
rect -960 280062 3575 280064
rect -960 279972 480 280062
rect 3509 280059 3575 280062
rect 555417 276450 555483 276453
rect 553380 276448 555483 276450
rect 553380 276392 555422 276448
rect 555478 276392 555483 276448
rect 553380 276390 555483 276392
rect 555417 276387 555483 276390
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 583520 272084 584960 272174
rect 8201 271826 8267 271829
rect 8201 271824 12052 271826
rect 8201 271768 8206 271824
rect 8262 271768 12052 271824
rect 8201 271766 12052 271768
rect 8201 271763 8267 271766
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 555417 264210 555483 264213
rect 553380 264208 555483 264210
rect 553380 264152 555422 264208
rect 555478 264152 555483 264208
rect 553380 264150 555483 264152
rect 555417 264147 555483 264150
rect 9397 259858 9463 259861
rect 9397 259856 12052 259858
rect 9397 259800 9402 259856
rect 9458 259800 12052 259856
rect 9397 259798 12052 259800
rect 9397 259795 9463 259798
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 556061 251970 556127 251973
rect 553380 251968 556127 251970
rect 553380 251912 556066 251968
rect 556122 251912 556127 251968
rect 553380 251910 556127 251912
rect 556061 251907 556127 251910
rect 8937 247890 9003 247893
rect 8937 247888 12052 247890
rect 8937 247832 8942 247888
rect 8998 247832 12052 247888
rect 8937 247830 12052 247832
rect 8937 247827 9003 247830
rect 579797 245578 579863 245581
rect 583520 245578 584960 245668
rect 579797 245576 584960 245578
rect 579797 245520 579802 245576
rect 579858 245520 584960 245576
rect 579797 245518 584960 245520
rect 579797 245515 579863 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3693 241090 3759 241093
rect -960 241088 3759 241090
rect -960 241032 3698 241088
rect 3754 241032 3759 241088
rect -960 241030 3759 241032
rect -960 240940 480 241030
rect 3693 241027 3759 241030
rect 555417 239730 555483 239733
rect 553380 239728 555483 239730
rect 553380 239672 555422 239728
rect 555478 239672 555483 239728
rect 553380 239670 555483 239672
rect 555417 239667 555483 239670
rect 9397 235922 9463 235925
rect 9397 235920 12052 235922
rect 9397 235864 9402 235920
rect 9458 235864 12052 235920
rect 9397 235862 12052 235864
rect 9397 235859 9463 235862
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 228034 480 228124
rect 4061 228034 4127 228037
rect -960 228032 4127 228034
rect -960 227976 4066 228032
rect 4122 227976 4127 228032
rect -960 227974 4127 227976
rect -960 227884 480 227974
rect 4061 227971 4127 227974
rect 555417 227490 555483 227493
rect 553380 227488 555483 227490
rect 553380 227432 555422 227488
rect 555478 227432 555483 227488
rect 553380 227430 555483 227432
rect 555417 227427 555483 227430
rect 8845 223954 8911 223957
rect 8845 223952 12052 223954
rect 8845 223896 8850 223952
rect 8906 223896 12052 223952
rect 8845 223894 12052 223896
rect 8845 223891 8911 223894
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 555417 215250 555483 215253
rect 553380 215248 555483 215250
rect 553380 215192 555422 215248
rect 555478 215192 555483 215248
rect 553380 215190 555483 215192
rect 555417 215187 555483 215190
rect -960 214978 480 215068
rect 3141 214978 3207 214981
rect -960 214976 3207 214978
rect -960 214920 3146 214976
rect 3202 214920 3207 214976
rect -960 214918 3207 214920
rect -960 214828 480 214918
rect 3141 214915 3207 214918
rect 9213 211986 9279 211989
rect 9213 211984 12052 211986
rect 9213 211928 9218 211984
rect 9274 211928 12052 211984
rect 9213 211926 12052 211928
rect 9213 211923 9279 211926
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 555417 203010 555483 203013
rect 553380 203008 555483 203010
rect 553380 202952 555422 203008
rect 555478 202952 555483 203008
rect 553380 202950 555483 202952
rect 555417 202947 555483 202950
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 8293 200018 8359 200021
rect 8293 200016 12052 200018
rect 8293 199960 8298 200016
rect 8354 199960 12052 200016
rect 8293 199958 12052 199960
rect 8293 199955 8359 199958
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 555417 190770 555483 190773
rect 553380 190768 555483 190770
rect 553380 190712 555422 190768
rect 555478 190712 555483 190768
rect 553380 190710 555483 190712
rect 555417 190707 555483 190710
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 9397 188050 9463 188053
rect 9397 188048 12052 188050
rect 9397 187992 9402 188048
rect 9458 187992 12052 188048
rect 9397 187990 12052 187992
rect 9397 187987 9463 187990
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 555417 178530 555483 178533
rect 553380 178528 555483 178530
rect 553380 178472 555422 178528
rect 555478 178472 555483 178528
rect 553380 178470 555483 178472
rect 555417 178467 555483 178470
rect 9397 176082 9463 176085
rect 9397 176080 12052 176082
rect -960 175946 480 176036
rect 9397 176024 9402 176080
rect 9458 176024 12052 176080
rect 9397 176022 12052 176024
rect 9397 176019 9463 176022
rect 3325 175946 3391 175949
rect -960 175944 3391 175946
rect -960 175888 3330 175944
rect 3386 175888 3391 175944
rect -960 175886 3391 175888
rect -960 175796 480 175886
rect 3325 175883 3391 175886
rect 555877 166290 555943 166293
rect 553380 166288 555943 166290
rect 553380 166232 555882 166288
rect 555938 166232 555943 166288
rect 553380 166230 555943 166232
rect 555877 166227 555943 166230
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 9397 164114 9463 164117
rect 9397 164112 12052 164114
rect 9397 164056 9402 164112
rect 9458 164056 12052 164112
rect 9397 164054 12052 164056
rect 9397 164051 9463 164054
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 555417 154050 555483 154053
rect 553380 154048 555483 154050
rect 553380 153992 555422 154048
rect 555478 153992 555483 154048
rect 553380 153990 555483 153992
rect 555417 153987 555483 153990
rect 579521 152690 579587 152693
rect 583520 152690 584960 152780
rect 579521 152688 584960 152690
rect 579521 152632 579526 152688
rect 579582 152632 584960 152688
rect 579521 152630 584960 152632
rect 579521 152627 579587 152630
rect 583520 152540 584960 152630
rect 8201 152146 8267 152149
rect 8201 152144 12052 152146
rect 8201 152088 8206 152144
rect 8262 152088 12052 152144
rect 8201 152086 12052 152088
rect 8201 152083 8267 152086
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 555417 141810 555483 141813
rect 553380 141808 555483 141810
rect 553380 141752 555422 141808
rect 555478 141752 555483 141808
rect 553380 141750 555483 141752
rect 555417 141747 555483 141750
rect 8201 140178 8267 140181
rect 8201 140176 12052 140178
rect 8201 140120 8206 140176
rect 8262 140120 12052 140176
rect 8201 140118 12052 140120
rect 8201 140115 8267 140118
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 555417 129570 555483 129573
rect 553380 129568 555483 129570
rect 553380 129512 555422 129568
rect 555478 129512 555483 129568
rect 553380 129510 555483 129512
rect 555417 129507 555483 129510
rect 8201 128210 8267 128213
rect 8201 128208 12052 128210
rect 8201 128152 8206 128208
rect 8262 128152 12052 128208
rect 8201 128150 12052 128152
rect 8201 128147 8267 128150
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 3417 123722 3483 123725
rect -960 123720 3483 123722
rect -960 123664 3422 123720
rect 3478 123664 3483 123720
rect -960 123662 3483 123664
rect -960 123572 480 123662
rect 3417 123659 3483 123662
rect 555417 117330 555483 117333
rect 553380 117328 555483 117330
rect 553380 117272 555422 117328
rect 555478 117272 555483 117328
rect 553380 117270 555483 117272
rect 555417 117267 555483 117270
rect 8937 116242 9003 116245
rect 8937 116240 12052 116242
rect 8937 116184 8942 116240
rect 8998 116184 12052 116240
rect 8937 116182 12052 116184
rect 8937 116179 9003 116182
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 555693 105090 555759 105093
rect 553380 105088 555759 105090
rect 553380 105032 555698 105088
rect 555754 105032 555759 105088
rect 553380 105030 555759 105032
rect 555693 105027 555759 105030
rect 9397 104274 9463 104277
rect 9397 104272 12052 104274
rect 9397 104216 9402 104272
rect 9458 104216 12052 104272
rect 9397 104214 12052 104216
rect 9397 104211 9463 104214
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 4061 97610 4127 97613
rect -960 97608 4127 97610
rect -960 97552 4066 97608
rect 4122 97552 4127 97608
rect -960 97550 4127 97552
rect -960 97460 480 97550
rect 4061 97547 4127 97550
rect 554773 92850 554839 92853
rect 553380 92848 554839 92850
rect 553380 92792 554778 92848
rect 554834 92792 554839 92848
rect 553380 92790 554839 92792
rect 554773 92787 554839 92790
rect 9397 92306 9463 92309
rect 9397 92304 12052 92306
rect 9397 92248 9402 92304
rect 9458 92248 12052 92304
rect 9397 92246 12052 92248
rect 9397 92243 9463 92246
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 4061 84690 4127 84693
rect -960 84688 4127 84690
rect -960 84632 4066 84688
rect 4122 84632 4127 84688
rect -960 84630 4127 84632
rect -960 84540 480 84630
rect 4061 84627 4127 84630
rect 555417 80610 555483 80613
rect 553380 80608 555483 80610
rect 553380 80552 555422 80608
rect 555478 80552 555483 80608
rect 553380 80550 555483 80552
rect 555417 80547 555483 80550
rect 8937 80338 9003 80341
rect 8937 80336 12052 80338
rect 8937 80280 8942 80336
rect 8998 80280 12052 80336
rect 8937 80278 12052 80280
rect 8937 80275 9003 80278
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 8937 68370 9003 68373
rect 555417 68370 555483 68373
rect 8937 68368 12052 68370
rect 8937 68312 8942 68368
rect 8998 68312 12052 68368
rect 8937 68310 12052 68312
rect 553380 68368 555483 68370
rect 553380 68312 555422 68368
rect 555478 68312 555483 68368
rect 553380 68310 555483 68312
rect 8937 68307 9003 68310
rect 555417 68307 555483 68310
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3141 58578 3207 58581
rect -960 58576 3207 58578
rect -960 58520 3146 58576
rect 3202 58520 3207 58576
rect -960 58518 3207 58520
rect -960 58428 480 58518
rect 3141 58515 3207 58518
rect 9397 56402 9463 56405
rect 9397 56400 12052 56402
rect 9397 56344 9402 56400
rect 9458 56344 12052 56400
rect 9397 56342 12052 56344
rect 9397 56339 9463 56342
rect 555417 56130 555483 56133
rect 553380 56128 555483 56130
rect 553380 56072 555422 56128
rect 555478 56072 555483 56128
rect 553380 56070 555483 56072
rect 555417 56067 555483 56070
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2773 45522 2839 45525
rect -960 45520 2839 45522
rect -960 45464 2778 45520
rect 2834 45464 2839 45520
rect -960 45462 2839 45464
rect -960 45372 480 45462
rect 2773 45459 2839 45462
rect 9397 44434 9463 44437
rect 9397 44432 12052 44434
rect 9397 44376 9402 44432
rect 9458 44376 12052 44432
rect 9397 44374 12052 44376
rect 9397 44371 9463 44374
rect 555417 43890 555483 43893
rect 553380 43888 555483 43890
rect 553380 43832 555422 43888
rect 555478 43832 555483 43888
rect 553380 43830 555483 43832
rect 555417 43827 555483 43830
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 9397 32466 9463 32469
rect 9397 32464 12052 32466
rect 9397 32408 9402 32464
rect 9458 32408 12052 32464
rect 9397 32406 12052 32408
rect 9397 32403 9463 32406
rect 555509 31650 555575 31653
rect 553380 31648 555575 31650
rect 553380 31592 555514 31648
rect 555570 31592 555575 31648
rect 553380 31590 555575 31592
rect 555509 31587 555575 31590
rect 9397 20498 9463 20501
rect 9397 20496 12052 20498
rect 9397 20440 9402 20496
rect 9458 20440 12052 20496
rect 9397 20438 12052 20440
rect 9397 20435 9463 20438
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect 555417 19410 555483 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect 553380 19408 555483 19410
rect 553380 19352 555422 19408
rect 555478 19352 555483 19408
rect 553380 19350 555483 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 555417 19347 555483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3141 6490 3207 6493
rect -960 6488 3207 6490
rect -960 6432 3146 6488
rect 3202 6432 3207 6488
rect 583520 6476 584960 6566
rect -960 6430 3207 6432
rect -960 6340 480 6430
rect 3141 6427 3207 6430
rect 39573 3362 39639 3365
rect 66253 3362 66319 3365
rect 39573 3360 66319 3362
rect 39573 3304 39578 3360
rect 39634 3304 66258 3360
rect 66314 3304 66319 3360
rect 39573 3302 66319 3304
rect 39573 3299 39639 3302
rect 66253 3299 66319 3302
rect 78581 3362 78647 3365
rect 99741 3362 99807 3365
rect 78581 3360 99807 3362
rect 78581 3304 78586 3360
rect 78642 3304 99746 3360
rect 99802 3304 99807 3360
rect 78581 3302 99807 3304
rect 78581 3299 78647 3302
rect 99741 3299 99807 3302
rect 458173 3362 458239 3365
rect 497089 3362 497155 3365
rect 458173 3360 497155 3362
rect 458173 3304 458178 3360
rect 458234 3304 497094 3360
rect 497150 3304 497155 3360
rect 458173 3302 497155 3304
rect 458173 3299 458239 3302
rect 497089 3299 497155 3302
rect 530025 3362 530091 3365
rect 582189 3362 582255 3365
rect 530025 3360 582255 3362
rect 530025 3304 530030 3360
rect 530086 3304 582194 3360
rect 582250 3304 582255 3360
rect 530025 3302 582255 3304
rect 530025 3299 530091 3302
rect 582189 3299 582255 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 660161 13574 662058
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 660161 17294 665778
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 660161 21014 669498
rect 24114 710598 24734 711590
rect 24114 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 24734 710598
rect 24114 710278 24734 710362
rect 24114 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 24734 710278
rect 24114 673774 24734 710042
rect 24114 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 24734 673774
rect 24114 673454 24734 673538
rect 24114 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 24734 673454
rect 24114 660161 24734 673218
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 27834 660161 28454 676938
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 660161 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 660161 42134 690618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 660161 45854 694338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 660161 49574 662058
rect 52674 708678 53294 711590
rect 52674 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 53294 708678
rect 52674 708358 53294 708442
rect 52674 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 53294 708358
rect 52674 666334 53294 708122
rect 52674 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 53294 666334
rect 52674 666014 53294 666098
rect 52674 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 53294 666014
rect 52674 660161 53294 665778
rect 56394 709638 57014 711590
rect 56394 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 57014 709638
rect 56394 709318 57014 709402
rect 56394 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 57014 709318
rect 56394 670054 57014 709082
rect 56394 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 57014 670054
rect 56394 669734 57014 669818
rect 56394 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 57014 669734
rect 56394 660161 57014 669498
rect 60114 710598 60734 711590
rect 60114 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 60734 710598
rect 60114 710278 60734 710362
rect 60114 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 60734 710278
rect 60114 673774 60734 710042
rect 60114 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 60734 673774
rect 60114 673454 60734 673538
rect 60114 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 60734 673454
rect 60114 660161 60734 673218
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 660161 64454 676938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 660161 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 663100 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 660161 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 660161 85574 662058
rect 88674 708678 89294 711590
rect 88674 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 89294 708678
rect 88674 708358 89294 708442
rect 88674 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 89294 708358
rect 88674 666334 89294 708122
rect 88674 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 89294 666334
rect 88674 666014 89294 666098
rect 88674 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 89294 666014
rect 88674 660161 89294 665778
rect 92394 709638 93014 711590
rect 92394 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 93014 709638
rect 92394 709318 93014 709402
rect 92394 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 93014 709318
rect 92394 670054 93014 709082
rect 92394 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 93014 670054
rect 92394 669734 93014 669818
rect 92394 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 93014 669734
rect 92394 663100 93014 669498
rect 96114 710598 96734 711590
rect 96114 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 96734 710598
rect 96114 710278 96734 710362
rect 96114 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 96734 710278
rect 96114 673774 96734 710042
rect 96114 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 96734 673774
rect 96114 673454 96734 673538
rect 96114 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 96734 673454
rect 96114 660161 96734 673218
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 660161 100454 676938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 660161 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 660161 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 660161 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 660161 121574 662058
rect 124674 708678 125294 711590
rect 124674 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 125294 708678
rect 124674 708358 125294 708442
rect 124674 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 125294 708358
rect 124674 666334 125294 708122
rect 124674 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 125294 666334
rect 124674 666014 125294 666098
rect 124674 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 125294 666014
rect 124674 660161 125294 665778
rect 128394 709638 129014 711590
rect 128394 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 129014 709638
rect 128394 709318 129014 709402
rect 128394 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 129014 709318
rect 128394 670054 129014 709082
rect 128394 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 129014 670054
rect 128394 669734 129014 669818
rect 128394 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 129014 669734
rect 128394 660161 129014 669498
rect 132114 710598 132734 711590
rect 132114 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 132734 710598
rect 132114 710278 132734 710362
rect 132114 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 132734 710278
rect 132114 673774 132734 710042
rect 132114 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 132734 673774
rect 132114 673454 132734 673538
rect 132114 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 132734 673454
rect 132114 660161 132734 673218
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 660161 136454 676938
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 660161 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 660161 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 660161 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 660161 157574 662058
rect 160674 708678 161294 711590
rect 160674 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 161294 708678
rect 160674 708358 161294 708442
rect 160674 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 161294 708358
rect 160674 666334 161294 708122
rect 160674 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 161294 666334
rect 160674 666014 161294 666098
rect 160674 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 161294 666014
rect 160674 660161 161294 665778
rect 164394 709638 165014 711590
rect 164394 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 165014 709638
rect 164394 709318 165014 709402
rect 164394 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 165014 709318
rect 164394 670054 165014 709082
rect 164394 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 165014 670054
rect 164394 669734 165014 669818
rect 164394 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 165014 669734
rect 164394 660161 165014 669498
rect 168114 710598 168734 711590
rect 168114 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 168734 710598
rect 168114 710278 168734 710362
rect 168114 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 168734 710278
rect 168114 673774 168734 710042
rect 168114 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 168734 673774
rect 168114 673454 168734 673538
rect 168114 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 168734 673454
rect 168114 660161 168734 673218
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 660161 172454 676938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 660161 182414 686898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 663100 186134 690618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 660161 189854 694338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 660161 193574 662058
rect 196674 708678 197294 711590
rect 196674 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 197294 708678
rect 196674 708358 197294 708442
rect 196674 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 197294 708358
rect 196674 666334 197294 708122
rect 196674 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 197294 666334
rect 196674 666014 197294 666098
rect 196674 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 197294 666014
rect 196674 660161 197294 665778
rect 200394 709638 201014 711590
rect 200394 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 201014 709638
rect 200394 709318 201014 709402
rect 200394 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 201014 709318
rect 200394 670054 201014 709082
rect 200394 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 201014 670054
rect 200394 669734 201014 669818
rect 200394 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 201014 669734
rect 200394 663100 201014 669498
rect 204114 710598 204734 711590
rect 204114 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 204734 710598
rect 204114 710278 204734 710362
rect 204114 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 204734 710278
rect 204114 673774 204734 710042
rect 204114 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 204734 673774
rect 204114 673454 204734 673538
rect 204114 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 204734 673454
rect 204114 660161 204734 673218
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 660161 208454 676938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 660161 218414 686898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 660161 222134 690618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 660161 225854 694338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 660161 229574 662058
rect 232674 708678 233294 711590
rect 232674 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 233294 708678
rect 232674 708358 233294 708442
rect 232674 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 233294 708358
rect 232674 666334 233294 708122
rect 232674 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 233294 666334
rect 232674 666014 233294 666098
rect 232674 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 233294 666014
rect 232674 660161 233294 665778
rect 236394 709638 237014 711590
rect 236394 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 237014 709638
rect 236394 709318 237014 709402
rect 236394 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 237014 709318
rect 236394 670054 237014 709082
rect 236394 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 237014 670054
rect 236394 669734 237014 669818
rect 236394 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 237014 669734
rect 236394 660161 237014 669498
rect 240114 710598 240734 711590
rect 240114 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 240734 710598
rect 240114 710278 240734 710362
rect 240114 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 240734 710278
rect 240114 673774 240734 710042
rect 240114 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 240734 673774
rect 240114 673454 240734 673538
rect 240114 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 240734 673454
rect 240114 660161 240734 673218
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 660161 244454 676938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 660161 254414 686898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 660161 258134 690618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 660161 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 660161 265574 662058
rect 268674 708678 269294 711590
rect 268674 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 269294 708678
rect 268674 708358 269294 708442
rect 268674 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 269294 708358
rect 268674 666334 269294 708122
rect 268674 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 269294 666334
rect 268674 666014 269294 666098
rect 268674 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 269294 666014
rect 268674 660161 269294 665778
rect 272394 709638 273014 711590
rect 272394 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 273014 709638
rect 272394 709318 273014 709402
rect 272394 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 273014 709318
rect 272394 670054 273014 709082
rect 272394 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 273014 670054
rect 272394 669734 273014 669818
rect 272394 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 273014 669734
rect 272394 660161 273014 669498
rect 276114 710598 276734 711590
rect 276114 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 276734 710598
rect 276114 710278 276734 710362
rect 276114 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 276734 710278
rect 276114 673774 276734 710042
rect 276114 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 276734 673774
rect 276114 673454 276734 673538
rect 276114 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 276734 673454
rect 276114 660161 276734 673218
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 660161 280454 676938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 660161 290414 686898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 660161 294134 690618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 660161 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 660161 301574 662058
rect 304674 708678 305294 711590
rect 304674 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 305294 708678
rect 304674 708358 305294 708442
rect 304674 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 305294 708358
rect 304674 666334 305294 708122
rect 304674 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 305294 666334
rect 304674 666014 305294 666098
rect 304674 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 305294 666014
rect 304674 660161 305294 665778
rect 308394 709638 309014 711590
rect 308394 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 309014 709638
rect 308394 709318 309014 709402
rect 308394 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 309014 709318
rect 308394 670054 309014 709082
rect 308394 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 309014 670054
rect 308394 669734 309014 669818
rect 308394 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 309014 669734
rect 308394 663100 309014 669498
rect 312114 710598 312734 711590
rect 312114 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 312734 710598
rect 312114 710278 312734 710362
rect 312114 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 312734 710278
rect 312114 673774 312734 710042
rect 312114 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 312734 673774
rect 312114 673454 312734 673538
rect 312114 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 312734 673454
rect 312114 660161 312734 673218
rect 315834 711558 316454 711590
rect 315834 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 316454 711558
rect 315834 711238 316454 711322
rect 315834 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 316454 711238
rect 315834 677494 316454 711002
rect 315834 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 316454 677494
rect 315834 677174 316454 677258
rect 315834 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 316454 677174
rect 315834 660161 316454 676938
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 660161 326414 686898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 660161 330134 690618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 660161 333854 694338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 660161 337574 662058
rect 340674 708678 341294 711590
rect 340674 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 341294 708678
rect 340674 708358 341294 708442
rect 340674 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 341294 708358
rect 340674 666334 341294 708122
rect 340674 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 341294 666334
rect 340674 666014 341294 666098
rect 340674 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 341294 666014
rect 340674 660161 341294 665778
rect 344394 709638 345014 711590
rect 344394 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 345014 709638
rect 344394 709318 345014 709402
rect 344394 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 345014 709318
rect 344394 670054 345014 709082
rect 344394 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 345014 670054
rect 344394 669734 345014 669818
rect 344394 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 345014 669734
rect 344394 660161 345014 669498
rect 348114 710598 348734 711590
rect 348114 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 348734 710598
rect 348114 710278 348734 710362
rect 348114 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 348734 710278
rect 348114 673774 348734 710042
rect 348114 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 348734 673774
rect 348114 673454 348734 673538
rect 348114 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 348734 673454
rect 348114 660161 348734 673218
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 660161 352454 676938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 660161 362414 686898
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 660161 366134 690618
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 663100 369854 694338
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 660161 373574 662058
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 660161 377294 665778
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 660161 381014 669498
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 660161 384734 673218
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 660161 388454 676938
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 660161 398414 686898
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 660161 402134 690618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 660161 405854 694338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 660161 409574 662058
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 660161 413294 665778
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 660161 417014 669498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 660161 420734 673218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 660161 424454 676938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 660161 434414 686898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 660161 438134 690618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 660161 441854 694338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 660161 445574 662058
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 448674 666334 449294 708122
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 660161 449294 665778
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 660161 453014 669498
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 660161 456734 673218
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 660161 460454 676938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 660161 470414 686898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 660161 474134 690618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 663100 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 660161 481574 662058
rect 484674 708678 485294 711590
rect 484674 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 485294 708678
rect 484674 708358 485294 708442
rect 484674 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 485294 708358
rect 484674 666334 485294 708122
rect 484674 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 485294 666334
rect 484674 666014 485294 666098
rect 484674 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 485294 666014
rect 484674 660161 485294 665778
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 660161 489014 669498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 663100 492734 673218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 660161 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 660161 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 660161 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 660161 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 660161 517574 662058
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 520674 660161 521294 665778
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 660161 525014 669498
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 528114 673774 528734 710042
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 660161 528734 673218
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 660161 532454 676938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 660161 542414 686898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 660161 546134 690618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 660161 549854 694338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 660161 553574 662058
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 31568 655174 31888 655206
rect 31568 654938 31610 655174
rect 31846 654938 31888 655174
rect 31568 654854 31888 654938
rect 31568 654618 31610 654854
rect 31846 654618 31888 654854
rect 31568 654586 31888 654618
rect 62288 655174 62608 655206
rect 62288 654938 62330 655174
rect 62566 654938 62608 655174
rect 62288 654854 62608 654938
rect 62288 654618 62330 654854
rect 62566 654618 62608 654854
rect 62288 654586 62608 654618
rect 93008 655174 93328 655206
rect 93008 654938 93050 655174
rect 93286 654938 93328 655174
rect 93008 654854 93328 654938
rect 93008 654618 93050 654854
rect 93286 654618 93328 654854
rect 93008 654586 93328 654618
rect 123728 655174 124048 655206
rect 123728 654938 123770 655174
rect 124006 654938 124048 655174
rect 123728 654854 124048 654938
rect 123728 654618 123770 654854
rect 124006 654618 124048 654854
rect 123728 654586 124048 654618
rect 154448 655174 154768 655206
rect 154448 654938 154490 655174
rect 154726 654938 154768 655174
rect 154448 654854 154768 654938
rect 154448 654618 154490 654854
rect 154726 654618 154768 654854
rect 154448 654586 154768 654618
rect 185168 655174 185488 655206
rect 185168 654938 185210 655174
rect 185446 654938 185488 655174
rect 185168 654854 185488 654938
rect 185168 654618 185210 654854
rect 185446 654618 185488 654854
rect 185168 654586 185488 654618
rect 215888 655174 216208 655206
rect 215888 654938 215930 655174
rect 216166 654938 216208 655174
rect 215888 654854 216208 654938
rect 215888 654618 215930 654854
rect 216166 654618 216208 654854
rect 215888 654586 216208 654618
rect 246608 655174 246928 655206
rect 246608 654938 246650 655174
rect 246886 654938 246928 655174
rect 246608 654854 246928 654938
rect 246608 654618 246650 654854
rect 246886 654618 246928 654854
rect 246608 654586 246928 654618
rect 277328 655174 277648 655206
rect 277328 654938 277370 655174
rect 277606 654938 277648 655174
rect 277328 654854 277648 654938
rect 277328 654618 277370 654854
rect 277606 654618 277648 654854
rect 277328 654586 277648 654618
rect 308048 655174 308368 655206
rect 308048 654938 308090 655174
rect 308326 654938 308368 655174
rect 308048 654854 308368 654938
rect 308048 654618 308090 654854
rect 308326 654618 308368 654854
rect 308048 654586 308368 654618
rect 338768 655174 339088 655206
rect 338768 654938 338810 655174
rect 339046 654938 339088 655174
rect 338768 654854 339088 654938
rect 338768 654618 338810 654854
rect 339046 654618 339088 654854
rect 338768 654586 339088 654618
rect 369488 655174 369808 655206
rect 369488 654938 369530 655174
rect 369766 654938 369808 655174
rect 369488 654854 369808 654938
rect 369488 654618 369530 654854
rect 369766 654618 369808 654854
rect 369488 654586 369808 654618
rect 400208 655174 400528 655206
rect 400208 654938 400250 655174
rect 400486 654938 400528 655174
rect 400208 654854 400528 654938
rect 400208 654618 400250 654854
rect 400486 654618 400528 654854
rect 400208 654586 400528 654618
rect 430928 655174 431248 655206
rect 430928 654938 430970 655174
rect 431206 654938 431248 655174
rect 430928 654854 431248 654938
rect 430928 654618 430970 654854
rect 431206 654618 431248 654854
rect 430928 654586 431248 654618
rect 461648 655174 461968 655206
rect 461648 654938 461690 655174
rect 461926 654938 461968 655174
rect 461648 654854 461968 654938
rect 461648 654618 461690 654854
rect 461926 654618 461968 654854
rect 461648 654586 461968 654618
rect 492368 655174 492688 655206
rect 492368 654938 492410 655174
rect 492646 654938 492688 655174
rect 492368 654854 492688 654938
rect 492368 654618 492410 654854
rect 492646 654618 492688 654854
rect 492368 654586 492688 654618
rect 523088 655174 523408 655206
rect 523088 654938 523130 655174
rect 523366 654938 523408 655174
rect 523088 654854 523408 654938
rect 523088 654618 523130 654854
rect 523366 654618 523408 654854
rect 523088 654586 523408 654618
rect 16208 651454 16528 651486
rect 16208 651218 16250 651454
rect 16486 651218 16528 651454
rect 16208 651134 16528 651218
rect 16208 650898 16250 651134
rect 16486 650898 16528 651134
rect 16208 650866 16528 650898
rect 46928 651454 47248 651486
rect 46928 651218 46970 651454
rect 47206 651218 47248 651454
rect 46928 651134 47248 651218
rect 46928 650898 46970 651134
rect 47206 650898 47248 651134
rect 46928 650866 47248 650898
rect 77648 651454 77968 651486
rect 77648 651218 77690 651454
rect 77926 651218 77968 651454
rect 77648 651134 77968 651218
rect 77648 650898 77690 651134
rect 77926 650898 77968 651134
rect 77648 650866 77968 650898
rect 108368 651454 108688 651486
rect 108368 651218 108410 651454
rect 108646 651218 108688 651454
rect 108368 651134 108688 651218
rect 108368 650898 108410 651134
rect 108646 650898 108688 651134
rect 108368 650866 108688 650898
rect 139088 651454 139408 651486
rect 139088 651218 139130 651454
rect 139366 651218 139408 651454
rect 139088 651134 139408 651218
rect 139088 650898 139130 651134
rect 139366 650898 139408 651134
rect 139088 650866 139408 650898
rect 169808 651454 170128 651486
rect 169808 651218 169850 651454
rect 170086 651218 170128 651454
rect 169808 651134 170128 651218
rect 169808 650898 169850 651134
rect 170086 650898 170128 651134
rect 169808 650866 170128 650898
rect 200528 651454 200848 651486
rect 200528 651218 200570 651454
rect 200806 651218 200848 651454
rect 200528 651134 200848 651218
rect 200528 650898 200570 651134
rect 200806 650898 200848 651134
rect 200528 650866 200848 650898
rect 231248 651454 231568 651486
rect 231248 651218 231290 651454
rect 231526 651218 231568 651454
rect 231248 651134 231568 651218
rect 231248 650898 231290 651134
rect 231526 650898 231568 651134
rect 231248 650866 231568 650898
rect 261968 651454 262288 651486
rect 261968 651218 262010 651454
rect 262246 651218 262288 651454
rect 261968 651134 262288 651218
rect 261968 650898 262010 651134
rect 262246 650898 262288 651134
rect 261968 650866 262288 650898
rect 292688 651454 293008 651486
rect 292688 651218 292730 651454
rect 292966 651218 293008 651454
rect 292688 651134 293008 651218
rect 292688 650898 292730 651134
rect 292966 650898 293008 651134
rect 292688 650866 293008 650898
rect 323408 651454 323728 651486
rect 323408 651218 323450 651454
rect 323686 651218 323728 651454
rect 323408 651134 323728 651218
rect 323408 650898 323450 651134
rect 323686 650898 323728 651134
rect 323408 650866 323728 650898
rect 354128 651454 354448 651486
rect 354128 651218 354170 651454
rect 354406 651218 354448 651454
rect 354128 651134 354448 651218
rect 354128 650898 354170 651134
rect 354406 650898 354448 651134
rect 354128 650866 354448 650898
rect 384848 651454 385168 651486
rect 384848 651218 384890 651454
rect 385126 651218 385168 651454
rect 384848 651134 385168 651218
rect 384848 650898 384890 651134
rect 385126 650898 385168 651134
rect 384848 650866 385168 650898
rect 415568 651454 415888 651486
rect 415568 651218 415610 651454
rect 415846 651218 415888 651454
rect 415568 651134 415888 651218
rect 415568 650898 415610 651134
rect 415846 650898 415888 651134
rect 415568 650866 415888 650898
rect 446288 651454 446608 651486
rect 446288 651218 446330 651454
rect 446566 651218 446608 651454
rect 446288 651134 446608 651218
rect 446288 650898 446330 651134
rect 446566 650898 446608 651134
rect 446288 650866 446608 650898
rect 477008 651454 477328 651486
rect 477008 651218 477050 651454
rect 477286 651218 477328 651454
rect 477008 651134 477328 651218
rect 477008 650898 477050 651134
rect 477286 650898 477328 651134
rect 477008 650866 477328 650898
rect 507728 651454 508048 651486
rect 507728 651218 507770 651454
rect 508006 651218 508048 651454
rect 507728 651134 508048 651218
rect 507728 650898 507770 651134
rect 508006 650898 508048 651134
rect 507728 650866 508048 650898
rect 538448 651454 538768 651486
rect 538448 651218 538490 651454
rect 538726 651218 538768 651454
rect 538448 651134 538768 651218
rect 538448 650898 538490 651134
rect 538726 650898 538768 651134
rect 538448 650866 538768 650898
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 31568 619174 31888 619206
rect 31568 618938 31610 619174
rect 31846 618938 31888 619174
rect 31568 618854 31888 618938
rect 31568 618618 31610 618854
rect 31846 618618 31888 618854
rect 31568 618586 31888 618618
rect 62288 619174 62608 619206
rect 62288 618938 62330 619174
rect 62566 618938 62608 619174
rect 62288 618854 62608 618938
rect 62288 618618 62330 618854
rect 62566 618618 62608 618854
rect 62288 618586 62608 618618
rect 93008 619174 93328 619206
rect 93008 618938 93050 619174
rect 93286 618938 93328 619174
rect 93008 618854 93328 618938
rect 93008 618618 93050 618854
rect 93286 618618 93328 618854
rect 93008 618586 93328 618618
rect 123728 619174 124048 619206
rect 123728 618938 123770 619174
rect 124006 618938 124048 619174
rect 123728 618854 124048 618938
rect 123728 618618 123770 618854
rect 124006 618618 124048 618854
rect 123728 618586 124048 618618
rect 154448 619174 154768 619206
rect 154448 618938 154490 619174
rect 154726 618938 154768 619174
rect 154448 618854 154768 618938
rect 154448 618618 154490 618854
rect 154726 618618 154768 618854
rect 154448 618586 154768 618618
rect 185168 619174 185488 619206
rect 185168 618938 185210 619174
rect 185446 618938 185488 619174
rect 185168 618854 185488 618938
rect 185168 618618 185210 618854
rect 185446 618618 185488 618854
rect 185168 618586 185488 618618
rect 215888 619174 216208 619206
rect 215888 618938 215930 619174
rect 216166 618938 216208 619174
rect 215888 618854 216208 618938
rect 215888 618618 215930 618854
rect 216166 618618 216208 618854
rect 215888 618586 216208 618618
rect 246608 619174 246928 619206
rect 246608 618938 246650 619174
rect 246886 618938 246928 619174
rect 246608 618854 246928 618938
rect 246608 618618 246650 618854
rect 246886 618618 246928 618854
rect 246608 618586 246928 618618
rect 277328 619174 277648 619206
rect 277328 618938 277370 619174
rect 277606 618938 277648 619174
rect 277328 618854 277648 618938
rect 277328 618618 277370 618854
rect 277606 618618 277648 618854
rect 277328 618586 277648 618618
rect 308048 619174 308368 619206
rect 308048 618938 308090 619174
rect 308326 618938 308368 619174
rect 308048 618854 308368 618938
rect 308048 618618 308090 618854
rect 308326 618618 308368 618854
rect 308048 618586 308368 618618
rect 338768 619174 339088 619206
rect 338768 618938 338810 619174
rect 339046 618938 339088 619174
rect 338768 618854 339088 618938
rect 338768 618618 338810 618854
rect 339046 618618 339088 618854
rect 338768 618586 339088 618618
rect 369488 619174 369808 619206
rect 369488 618938 369530 619174
rect 369766 618938 369808 619174
rect 369488 618854 369808 618938
rect 369488 618618 369530 618854
rect 369766 618618 369808 618854
rect 369488 618586 369808 618618
rect 400208 619174 400528 619206
rect 400208 618938 400250 619174
rect 400486 618938 400528 619174
rect 400208 618854 400528 618938
rect 400208 618618 400250 618854
rect 400486 618618 400528 618854
rect 400208 618586 400528 618618
rect 430928 619174 431248 619206
rect 430928 618938 430970 619174
rect 431206 618938 431248 619174
rect 430928 618854 431248 618938
rect 430928 618618 430970 618854
rect 431206 618618 431248 618854
rect 430928 618586 431248 618618
rect 461648 619174 461968 619206
rect 461648 618938 461690 619174
rect 461926 618938 461968 619174
rect 461648 618854 461968 618938
rect 461648 618618 461690 618854
rect 461926 618618 461968 618854
rect 461648 618586 461968 618618
rect 492368 619174 492688 619206
rect 492368 618938 492410 619174
rect 492646 618938 492688 619174
rect 492368 618854 492688 618938
rect 492368 618618 492410 618854
rect 492646 618618 492688 618854
rect 492368 618586 492688 618618
rect 523088 619174 523408 619206
rect 523088 618938 523130 619174
rect 523366 618938 523408 619174
rect 523088 618854 523408 618938
rect 523088 618618 523130 618854
rect 523366 618618 523408 618854
rect 523088 618586 523408 618618
rect 16208 615454 16528 615486
rect 16208 615218 16250 615454
rect 16486 615218 16528 615454
rect 16208 615134 16528 615218
rect 16208 614898 16250 615134
rect 16486 614898 16528 615134
rect 16208 614866 16528 614898
rect 46928 615454 47248 615486
rect 46928 615218 46970 615454
rect 47206 615218 47248 615454
rect 46928 615134 47248 615218
rect 46928 614898 46970 615134
rect 47206 614898 47248 615134
rect 46928 614866 47248 614898
rect 77648 615454 77968 615486
rect 77648 615218 77690 615454
rect 77926 615218 77968 615454
rect 77648 615134 77968 615218
rect 77648 614898 77690 615134
rect 77926 614898 77968 615134
rect 77648 614866 77968 614898
rect 108368 615454 108688 615486
rect 108368 615218 108410 615454
rect 108646 615218 108688 615454
rect 108368 615134 108688 615218
rect 108368 614898 108410 615134
rect 108646 614898 108688 615134
rect 108368 614866 108688 614898
rect 139088 615454 139408 615486
rect 139088 615218 139130 615454
rect 139366 615218 139408 615454
rect 139088 615134 139408 615218
rect 139088 614898 139130 615134
rect 139366 614898 139408 615134
rect 139088 614866 139408 614898
rect 169808 615454 170128 615486
rect 169808 615218 169850 615454
rect 170086 615218 170128 615454
rect 169808 615134 170128 615218
rect 169808 614898 169850 615134
rect 170086 614898 170128 615134
rect 169808 614866 170128 614898
rect 200528 615454 200848 615486
rect 200528 615218 200570 615454
rect 200806 615218 200848 615454
rect 200528 615134 200848 615218
rect 200528 614898 200570 615134
rect 200806 614898 200848 615134
rect 200528 614866 200848 614898
rect 231248 615454 231568 615486
rect 231248 615218 231290 615454
rect 231526 615218 231568 615454
rect 231248 615134 231568 615218
rect 231248 614898 231290 615134
rect 231526 614898 231568 615134
rect 231248 614866 231568 614898
rect 261968 615454 262288 615486
rect 261968 615218 262010 615454
rect 262246 615218 262288 615454
rect 261968 615134 262288 615218
rect 261968 614898 262010 615134
rect 262246 614898 262288 615134
rect 261968 614866 262288 614898
rect 292688 615454 293008 615486
rect 292688 615218 292730 615454
rect 292966 615218 293008 615454
rect 292688 615134 293008 615218
rect 292688 614898 292730 615134
rect 292966 614898 293008 615134
rect 292688 614866 293008 614898
rect 323408 615454 323728 615486
rect 323408 615218 323450 615454
rect 323686 615218 323728 615454
rect 323408 615134 323728 615218
rect 323408 614898 323450 615134
rect 323686 614898 323728 615134
rect 323408 614866 323728 614898
rect 354128 615454 354448 615486
rect 354128 615218 354170 615454
rect 354406 615218 354448 615454
rect 354128 615134 354448 615218
rect 354128 614898 354170 615134
rect 354406 614898 354448 615134
rect 354128 614866 354448 614898
rect 384848 615454 385168 615486
rect 384848 615218 384890 615454
rect 385126 615218 385168 615454
rect 384848 615134 385168 615218
rect 384848 614898 384890 615134
rect 385126 614898 385168 615134
rect 384848 614866 385168 614898
rect 415568 615454 415888 615486
rect 415568 615218 415610 615454
rect 415846 615218 415888 615454
rect 415568 615134 415888 615218
rect 415568 614898 415610 615134
rect 415846 614898 415888 615134
rect 415568 614866 415888 614898
rect 446288 615454 446608 615486
rect 446288 615218 446330 615454
rect 446566 615218 446608 615454
rect 446288 615134 446608 615218
rect 446288 614898 446330 615134
rect 446566 614898 446608 615134
rect 446288 614866 446608 614898
rect 477008 615454 477328 615486
rect 477008 615218 477050 615454
rect 477286 615218 477328 615454
rect 477008 615134 477328 615218
rect 477008 614898 477050 615134
rect 477286 614898 477328 615134
rect 477008 614866 477328 614898
rect 507728 615454 508048 615486
rect 507728 615218 507770 615454
rect 508006 615218 508048 615454
rect 507728 615134 508048 615218
rect 507728 614898 507770 615134
rect 508006 614898 508048 615134
rect 507728 614866 508048 614898
rect 538448 615454 538768 615486
rect 538448 615218 538490 615454
rect 538726 615218 538768 615454
rect 538448 615134 538768 615218
rect 538448 614898 538490 615134
rect 538726 614898 538768 615134
rect 538448 614866 538768 614898
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 31568 583174 31888 583206
rect 31568 582938 31610 583174
rect 31846 582938 31888 583174
rect 31568 582854 31888 582938
rect 31568 582618 31610 582854
rect 31846 582618 31888 582854
rect 31568 582586 31888 582618
rect 62288 583174 62608 583206
rect 62288 582938 62330 583174
rect 62566 582938 62608 583174
rect 62288 582854 62608 582938
rect 62288 582618 62330 582854
rect 62566 582618 62608 582854
rect 62288 582586 62608 582618
rect 93008 583174 93328 583206
rect 93008 582938 93050 583174
rect 93286 582938 93328 583174
rect 93008 582854 93328 582938
rect 93008 582618 93050 582854
rect 93286 582618 93328 582854
rect 93008 582586 93328 582618
rect 123728 583174 124048 583206
rect 123728 582938 123770 583174
rect 124006 582938 124048 583174
rect 123728 582854 124048 582938
rect 123728 582618 123770 582854
rect 124006 582618 124048 582854
rect 123728 582586 124048 582618
rect 154448 583174 154768 583206
rect 154448 582938 154490 583174
rect 154726 582938 154768 583174
rect 154448 582854 154768 582938
rect 154448 582618 154490 582854
rect 154726 582618 154768 582854
rect 154448 582586 154768 582618
rect 185168 583174 185488 583206
rect 185168 582938 185210 583174
rect 185446 582938 185488 583174
rect 185168 582854 185488 582938
rect 185168 582618 185210 582854
rect 185446 582618 185488 582854
rect 185168 582586 185488 582618
rect 215888 583174 216208 583206
rect 215888 582938 215930 583174
rect 216166 582938 216208 583174
rect 215888 582854 216208 582938
rect 215888 582618 215930 582854
rect 216166 582618 216208 582854
rect 215888 582586 216208 582618
rect 246608 583174 246928 583206
rect 246608 582938 246650 583174
rect 246886 582938 246928 583174
rect 246608 582854 246928 582938
rect 246608 582618 246650 582854
rect 246886 582618 246928 582854
rect 246608 582586 246928 582618
rect 277328 583174 277648 583206
rect 277328 582938 277370 583174
rect 277606 582938 277648 583174
rect 277328 582854 277648 582938
rect 277328 582618 277370 582854
rect 277606 582618 277648 582854
rect 277328 582586 277648 582618
rect 308048 583174 308368 583206
rect 308048 582938 308090 583174
rect 308326 582938 308368 583174
rect 308048 582854 308368 582938
rect 308048 582618 308090 582854
rect 308326 582618 308368 582854
rect 308048 582586 308368 582618
rect 338768 583174 339088 583206
rect 338768 582938 338810 583174
rect 339046 582938 339088 583174
rect 338768 582854 339088 582938
rect 338768 582618 338810 582854
rect 339046 582618 339088 582854
rect 338768 582586 339088 582618
rect 369488 583174 369808 583206
rect 369488 582938 369530 583174
rect 369766 582938 369808 583174
rect 369488 582854 369808 582938
rect 369488 582618 369530 582854
rect 369766 582618 369808 582854
rect 369488 582586 369808 582618
rect 400208 583174 400528 583206
rect 400208 582938 400250 583174
rect 400486 582938 400528 583174
rect 400208 582854 400528 582938
rect 400208 582618 400250 582854
rect 400486 582618 400528 582854
rect 400208 582586 400528 582618
rect 430928 583174 431248 583206
rect 430928 582938 430970 583174
rect 431206 582938 431248 583174
rect 430928 582854 431248 582938
rect 430928 582618 430970 582854
rect 431206 582618 431248 582854
rect 430928 582586 431248 582618
rect 461648 583174 461968 583206
rect 461648 582938 461690 583174
rect 461926 582938 461968 583174
rect 461648 582854 461968 582938
rect 461648 582618 461690 582854
rect 461926 582618 461968 582854
rect 461648 582586 461968 582618
rect 492368 583174 492688 583206
rect 492368 582938 492410 583174
rect 492646 582938 492688 583174
rect 492368 582854 492688 582938
rect 492368 582618 492410 582854
rect 492646 582618 492688 582854
rect 492368 582586 492688 582618
rect 523088 583174 523408 583206
rect 523088 582938 523130 583174
rect 523366 582938 523408 583174
rect 523088 582854 523408 582938
rect 523088 582618 523130 582854
rect 523366 582618 523408 582854
rect 523088 582586 523408 582618
rect 16208 579454 16528 579486
rect 16208 579218 16250 579454
rect 16486 579218 16528 579454
rect 16208 579134 16528 579218
rect 16208 578898 16250 579134
rect 16486 578898 16528 579134
rect 16208 578866 16528 578898
rect 46928 579454 47248 579486
rect 46928 579218 46970 579454
rect 47206 579218 47248 579454
rect 46928 579134 47248 579218
rect 46928 578898 46970 579134
rect 47206 578898 47248 579134
rect 46928 578866 47248 578898
rect 77648 579454 77968 579486
rect 77648 579218 77690 579454
rect 77926 579218 77968 579454
rect 77648 579134 77968 579218
rect 77648 578898 77690 579134
rect 77926 578898 77968 579134
rect 77648 578866 77968 578898
rect 108368 579454 108688 579486
rect 108368 579218 108410 579454
rect 108646 579218 108688 579454
rect 108368 579134 108688 579218
rect 108368 578898 108410 579134
rect 108646 578898 108688 579134
rect 108368 578866 108688 578898
rect 139088 579454 139408 579486
rect 139088 579218 139130 579454
rect 139366 579218 139408 579454
rect 139088 579134 139408 579218
rect 139088 578898 139130 579134
rect 139366 578898 139408 579134
rect 139088 578866 139408 578898
rect 169808 579454 170128 579486
rect 169808 579218 169850 579454
rect 170086 579218 170128 579454
rect 169808 579134 170128 579218
rect 169808 578898 169850 579134
rect 170086 578898 170128 579134
rect 169808 578866 170128 578898
rect 200528 579454 200848 579486
rect 200528 579218 200570 579454
rect 200806 579218 200848 579454
rect 200528 579134 200848 579218
rect 200528 578898 200570 579134
rect 200806 578898 200848 579134
rect 200528 578866 200848 578898
rect 231248 579454 231568 579486
rect 231248 579218 231290 579454
rect 231526 579218 231568 579454
rect 231248 579134 231568 579218
rect 231248 578898 231290 579134
rect 231526 578898 231568 579134
rect 231248 578866 231568 578898
rect 261968 579454 262288 579486
rect 261968 579218 262010 579454
rect 262246 579218 262288 579454
rect 261968 579134 262288 579218
rect 261968 578898 262010 579134
rect 262246 578898 262288 579134
rect 261968 578866 262288 578898
rect 292688 579454 293008 579486
rect 292688 579218 292730 579454
rect 292966 579218 293008 579454
rect 292688 579134 293008 579218
rect 292688 578898 292730 579134
rect 292966 578898 293008 579134
rect 292688 578866 293008 578898
rect 323408 579454 323728 579486
rect 323408 579218 323450 579454
rect 323686 579218 323728 579454
rect 323408 579134 323728 579218
rect 323408 578898 323450 579134
rect 323686 578898 323728 579134
rect 323408 578866 323728 578898
rect 354128 579454 354448 579486
rect 354128 579218 354170 579454
rect 354406 579218 354448 579454
rect 354128 579134 354448 579218
rect 354128 578898 354170 579134
rect 354406 578898 354448 579134
rect 354128 578866 354448 578898
rect 384848 579454 385168 579486
rect 384848 579218 384890 579454
rect 385126 579218 385168 579454
rect 384848 579134 385168 579218
rect 384848 578898 384890 579134
rect 385126 578898 385168 579134
rect 384848 578866 385168 578898
rect 415568 579454 415888 579486
rect 415568 579218 415610 579454
rect 415846 579218 415888 579454
rect 415568 579134 415888 579218
rect 415568 578898 415610 579134
rect 415846 578898 415888 579134
rect 415568 578866 415888 578898
rect 446288 579454 446608 579486
rect 446288 579218 446330 579454
rect 446566 579218 446608 579454
rect 446288 579134 446608 579218
rect 446288 578898 446330 579134
rect 446566 578898 446608 579134
rect 446288 578866 446608 578898
rect 477008 579454 477328 579486
rect 477008 579218 477050 579454
rect 477286 579218 477328 579454
rect 477008 579134 477328 579218
rect 477008 578898 477050 579134
rect 477286 578898 477328 579134
rect 477008 578866 477328 578898
rect 507728 579454 508048 579486
rect 507728 579218 507770 579454
rect 508006 579218 508048 579454
rect 507728 579134 508048 579218
rect 507728 578898 507770 579134
rect 508006 578898 508048 579134
rect 507728 578866 508048 578898
rect 538448 579454 538768 579486
rect 538448 579218 538490 579454
rect 538726 579218 538768 579454
rect 538448 579134 538768 579218
rect 538448 578898 538490 579134
rect 538726 578898 538768 579134
rect 538448 578866 538768 578898
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 31568 547174 31888 547206
rect 31568 546938 31610 547174
rect 31846 546938 31888 547174
rect 31568 546854 31888 546938
rect 31568 546618 31610 546854
rect 31846 546618 31888 546854
rect 31568 546586 31888 546618
rect 62288 547174 62608 547206
rect 62288 546938 62330 547174
rect 62566 546938 62608 547174
rect 62288 546854 62608 546938
rect 62288 546618 62330 546854
rect 62566 546618 62608 546854
rect 62288 546586 62608 546618
rect 93008 547174 93328 547206
rect 93008 546938 93050 547174
rect 93286 546938 93328 547174
rect 93008 546854 93328 546938
rect 93008 546618 93050 546854
rect 93286 546618 93328 546854
rect 93008 546586 93328 546618
rect 123728 547174 124048 547206
rect 123728 546938 123770 547174
rect 124006 546938 124048 547174
rect 123728 546854 124048 546938
rect 123728 546618 123770 546854
rect 124006 546618 124048 546854
rect 123728 546586 124048 546618
rect 154448 547174 154768 547206
rect 154448 546938 154490 547174
rect 154726 546938 154768 547174
rect 154448 546854 154768 546938
rect 154448 546618 154490 546854
rect 154726 546618 154768 546854
rect 154448 546586 154768 546618
rect 185168 547174 185488 547206
rect 185168 546938 185210 547174
rect 185446 546938 185488 547174
rect 185168 546854 185488 546938
rect 185168 546618 185210 546854
rect 185446 546618 185488 546854
rect 185168 546586 185488 546618
rect 215888 547174 216208 547206
rect 215888 546938 215930 547174
rect 216166 546938 216208 547174
rect 215888 546854 216208 546938
rect 215888 546618 215930 546854
rect 216166 546618 216208 546854
rect 215888 546586 216208 546618
rect 246608 547174 246928 547206
rect 246608 546938 246650 547174
rect 246886 546938 246928 547174
rect 246608 546854 246928 546938
rect 246608 546618 246650 546854
rect 246886 546618 246928 546854
rect 246608 546586 246928 546618
rect 277328 547174 277648 547206
rect 277328 546938 277370 547174
rect 277606 546938 277648 547174
rect 277328 546854 277648 546938
rect 277328 546618 277370 546854
rect 277606 546618 277648 546854
rect 277328 546586 277648 546618
rect 308048 547174 308368 547206
rect 308048 546938 308090 547174
rect 308326 546938 308368 547174
rect 308048 546854 308368 546938
rect 308048 546618 308090 546854
rect 308326 546618 308368 546854
rect 308048 546586 308368 546618
rect 338768 547174 339088 547206
rect 338768 546938 338810 547174
rect 339046 546938 339088 547174
rect 338768 546854 339088 546938
rect 338768 546618 338810 546854
rect 339046 546618 339088 546854
rect 338768 546586 339088 546618
rect 369488 547174 369808 547206
rect 369488 546938 369530 547174
rect 369766 546938 369808 547174
rect 369488 546854 369808 546938
rect 369488 546618 369530 546854
rect 369766 546618 369808 546854
rect 369488 546586 369808 546618
rect 400208 547174 400528 547206
rect 400208 546938 400250 547174
rect 400486 546938 400528 547174
rect 400208 546854 400528 546938
rect 400208 546618 400250 546854
rect 400486 546618 400528 546854
rect 400208 546586 400528 546618
rect 430928 547174 431248 547206
rect 430928 546938 430970 547174
rect 431206 546938 431248 547174
rect 430928 546854 431248 546938
rect 430928 546618 430970 546854
rect 431206 546618 431248 546854
rect 430928 546586 431248 546618
rect 461648 547174 461968 547206
rect 461648 546938 461690 547174
rect 461926 546938 461968 547174
rect 461648 546854 461968 546938
rect 461648 546618 461690 546854
rect 461926 546618 461968 546854
rect 461648 546586 461968 546618
rect 492368 547174 492688 547206
rect 492368 546938 492410 547174
rect 492646 546938 492688 547174
rect 492368 546854 492688 546938
rect 492368 546618 492410 546854
rect 492646 546618 492688 546854
rect 492368 546586 492688 546618
rect 523088 547174 523408 547206
rect 523088 546938 523130 547174
rect 523366 546938 523408 547174
rect 523088 546854 523408 546938
rect 523088 546618 523130 546854
rect 523366 546618 523408 546854
rect 523088 546586 523408 546618
rect 16208 543454 16528 543486
rect 16208 543218 16250 543454
rect 16486 543218 16528 543454
rect 16208 543134 16528 543218
rect 16208 542898 16250 543134
rect 16486 542898 16528 543134
rect 16208 542866 16528 542898
rect 46928 543454 47248 543486
rect 46928 543218 46970 543454
rect 47206 543218 47248 543454
rect 46928 543134 47248 543218
rect 46928 542898 46970 543134
rect 47206 542898 47248 543134
rect 46928 542866 47248 542898
rect 77648 543454 77968 543486
rect 77648 543218 77690 543454
rect 77926 543218 77968 543454
rect 77648 543134 77968 543218
rect 77648 542898 77690 543134
rect 77926 542898 77968 543134
rect 77648 542866 77968 542898
rect 108368 543454 108688 543486
rect 108368 543218 108410 543454
rect 108646 543218 108688 543454
rect 108368 543134 108688 543218
rect 108368 542898 108410 543134
rect 108646 542898 108688 543134
rect 108368 542866 108688 542898
rect 139088 543454 139408 543486
rect 139088 543218 139130 543454
rect 139366 543218 139408 543454
rect 139088 543134 139408 543218
rect 139088 542898 139130 543134
rect 139366 542898 139408 543134
rect 139088 542866 139408 542898
rect 169808 543454 170128 543486
rect 169808 543218 169850 543454
rect 170086 543218 170128 543454
rect 169808 543134 170128 543218
rect 169808 542898 169850 543134
rect 170086 542898 170128 543134
rect 169808 542866 170128 542898
rect 200528 543454 200848 543486
rect 200528 543218 200570 543454
rect 200806 543218 200848 543454
rect 200528 543134 200848 543218
rect 200528 542898 200570 543134
rect 200806 542898 200848 543134
rect 200528 542866 200848 542898
rect 231248 543454 231568 543486
rect 231248 543218 231290 543454
rect 231526 543218 231568 543454
rect 231248 543134 231568 543218
rect 231248 542898 231290 543134
rect 231526 542898 231568 543134
rect 231248 542866 231568 542898
rect 261968 543454 262288 543486
rect 261968 543218 262010 543454
rect 262246 543218 262288 543454
rect 261968 543134 262288 543218
rect 261968 542898 262010 543134
rect 262246 542898 262288 543134
rect 261968 542866 262288 542898
rect 292688 543454 293008 543486
rect 292688 543218 292730 543454
rect 292966 543218 293008 543454
rect 292688 543134 293008 543218
rect 292688 542898 292730 543134
rect 292966 542898 293008 543134
rect 292688 542866 293008 542898
rect 323408 543454 323728 543486
rect 323408 543218 323450 543454
rect 323686 543218 323728 543454
rect 323408 543134 323728 543218
rect 323408 542898 323450 543134
rect 323686 542898 323728 543134
rect 323408 542866 323728 542898
rect 354128 543454 354448 543486
rect 354128 543218 354170 543454
rect 354406 543218 354448 543454
rect 354128 543134 354448 543218
rect 354128 542898 354170 543134
rect 354406 542898 354448 543134
rect 354128 542866 354448 542898
rect 384848 543454 385168 543486
rect 384848 543218 384890 543454
rect 385126 543218 385168 543454
rect 384848 543134 385168 543218
rect 384848 542898 384890 543134
rect 385126 542898 385168 543134
rect 384848 542866 385168 542898
rect 415568 543454 415888 543486
rect 415568 543218 415610 543454
rect 415846 543218 415888 543454
rect 415568 543134 415888 543218
rect 415568 542898 415610 543134
rect 415846 542898 415888 543134
rect 415568 542866 415888 542898
rect 446288 543454 446608 543486
rect 446288 543218 446330 543454
rect 446566 543218 446608 543454
rect 446288 543134 446608 543218
rect 446288 542898 446330 543134
rect 446566 542898 446608 543134
rect 446288 542866 446608 542898
rect 477008 543454 477328 543486
rect 477008 543218 477050 543454
rect 477286 543218 477328 543454
rect 477008 543134 477328 543218
rect 477008 542898 477050 543134
rect 477286 542898 477328 543134
rect 477008 542866 477328 542898
rect 507728 543454 508048 543486
rect 507728 543218 507770 543454
rect 508006 543218 508048 543454
rect 507728 543134 508048 543218
rect 507728 542898 507770 543134
rect 508006 542898 508048 543134
rect 507728 542866 508048 542898
rect 538448 543454 538768 543486
rect 538448 543218 538490 543454
rect 538726 543218 538768 543454
rect 538448 543134 538768 543218
rect 538448 542898 538490 543134
rect 538726 542898 538768 543134
rect 538448 542866 538768 542898
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 31568 511174 31888 511206
rect 31568 510938 31610 511174
rect 31846 510938 31888 511174
rect 31568 510854 31888 510938
rect 31568 510618 31610 510854
rect 31846 510618 31888 510854
rect 31568 510586 31888 510618
rect 62288 511174 62608 511206
rect 62288 510938 62330 511174
rect 62566 510938 62608 511174
rect 62288 510854 62608 510938
rect 62288 510618 62330 510854
rect 62566 510618 62608 510854
rect 62288 510586 62608 510618
rect 93008 511174 93328 511206
rect 93008 510938 93050 511174
rect 93286 510938 93328 511174
rect 93008 510854 93328 510938
rect 93008 510618 93050 510854
rect 93286 510618 93328 510854
rect 93008 510586 93328 510618
rect 123728 511174 124048 511206
rect 123728 510938 123770 511174
rect 124006 510938 124048 511174
rect 123728 510854 124048 510938
rect 123728 510618 123770 510854
rect 124006 510618 124048 510854
rect 123728 510586 124048 510618
rect 154448 511174 154768 511206
rect 154448 510938 154490 511174
rect 154726 510938 154768 511174
rect 154448 510854 154768 510938
rect 154448 510618 154490 510854
rect 154726 510618 154768 510854
rect 154448 510586 154768 510618
rect 185168 511174 185488 511206
rect 185168 510938 185210 511174
rect 185446 510938 185488 511174
rect 185168 510854 185488 510938
rect 185168 510618 185210 510854
rect 185446 510618 185488 510854
rect 185168 510586 185488 510618
rect 215888 511174 216208 511206
rect 215888 510938 215930 511174
rect 216166 510938 216208 511174
rect 215888 510854 216208 510938
rect 215888 510618 215930 510854
rect 216166 510618 216208 510854
rect 215888 510586 216208 510618
rect 246608 511174 246928 511206
rect 246608 510938 246650 511174
rect 246886 510938 246928 511174
rect 246608 510854 246928 510938
rect 246608 510618 246650 510854
rect 246886 510618 246928 510854
rect 246608 510586 246928 510618
rect 277328 511174 277648 511206
rect 277328 510938 277370 511174
rect 277606 510938 277648 511174
rect 277328 510854 277648 510938
rect 277328 510618 277370 510854
rect 277606 510618 277648 510854
rect 277328 510586 277648 510618
rect 308048 511174 308368 511206
rect 308048 510938 308090 511174
rect 308326 510938 308368 511174
rect 308048 510854 308368 510938
rect 308048 510618 308090 510854
rect 308326 510618 308368 510854
rect 308048 510586 308368 510618
rect 338768 511174 339088 511206
rect 338768 510938 338810 511174
rect 339046 510938 339088 511174
rect 338768 510854 339088 510938
rect 338768 510618 338810 510854
rect 339046 510618 339088 510854
rect 338768 510586 339088 510618
rect 369488 511174 369808 511206
rect 369488 510938 369530 511174
rect 369766 510938 369808 511174
rect 369488 510854 369808 510938
rect 369488 510618 369530 510854
rect 369766 510618 369808 510854
rect 369488 510586 369808 510618
rect 400208 511174 400528 511206
rect 400208 510938 400250 511174
rect 400486 510938 400528 511174
rect 400208 510854 400528 510938
rect 400208 510618 400250 510854
rect 400486 510618 400528 510854
rect 400208 510586 400528 510618
rect 430928 511174 431248 511206
rect 430928 510938 430970 511174
rect 431206 510938 431248 511174
rect 430928 510854 431248 510938
rect 430928 510618 430970 510854
rect 431206 510618 431248 510854
rect 430928 510586 431248 510618
rect 461648 511174 461968 511206
rect 461648 510938 461690 511174
rect 461926 510938 461968 511174
rect 461648 510854 461968 510938
rect 461648 510618 461690 510854
rect 461926 510618 461968 510854
rect 461648 510586 461968 510618
rect 492368 511174 492688 511206
rect 492368 510938 492410 511174
rect 492646 510938 492688 511174
rect 492368 510854 492688 510938
rect 492368 510618 492410 510854
rect 492646 510618 492688 510854
rect 492368 510586 492688 510618
rect 523088 511174 523408 511206
rect 523088 510938 523130 511174
rect 523366 510938 523408 511174
rect 523088 510854 523408 510938
rect 523088 510618 523130 510854
rect 523366 510618 523408 510854
rect 523088 510586 523408 510618
rect 16208 507454 16528 507486
rect 16208 507218 16250 507454
rect 16486 507218 16528 507454
rect 16208 507134 16528 507218
rect 16208 506898 16250 507134
rect 16486 506898 16528 507134
rect 16208 506866 16528 506898
rect 46928 507454 47248 507486
rect 46928 507218 46970 507454
rect 47206 507218 47248 507454
rect 46928 507134 47248 507218
rect 46928 506898 46970 507134
rect 47206 506898 47248 507134
rect 46928 506866 47248 506898
rect 77648 507454 77968 507486
rect 77648 507218 77690 507454
rect 77926 507218 77968 507454
rect 77648 507134 77968 507218
rect 77648 506898 77690 507134
rect 77926 506898 77968 507134
rect 77648 506866 77968 506898
rect 108368 507454 108688 507486
rect 108368 507218 108410 507454
rect 108646 507218 108688 507454
rect 108368 507134 108688 507218
rect 108368 506898 108410 507134
rect 108646 506898 108688 507134
rect 108368 506866 108688 506898
rect 139088 507454 139408 507486
rect 139088 507218 139130 507454
rect 139366 507218 139408 507454
rect 139088 507134 139408 507218
rect 139088 506898 139130 507134
rect 139366 506898 139408 507134
rect 139088 506866 139408 506898
rect 169808 507454 170128 507486
rect 169808 507218 169850 507454
rect 170086 507218 170128 507454
rect 169808 507134 170128 507218
rect 169808 506898 169850 507134
rect 170086 506898 170128 507134
rect 169808 506866 170128 506898
rect 200528 507454 200848 507486
rect 200528 507218 200570 507454
rect 200806 507218 200848 507454
rect 200528 507134 200848 507218
rect 200528 506898 200570 507134
rect 200806 506898 200848 507134
rect 200528 506866 200848 506898
rect 231248 507454 231568 507486
rect 231248 507218 231290 507454
rect 231526 507218 231568 507454
rect 231248 507134 231568 507218
rect 231248 506898 231290 507134
rect 231526 506898 231568 507134
rect 231248 506866 231568 506898
rect 261968 507454 262288 507486
rect 261968 507218 262010 507454
rect 262246 507218 262288 507454
rect 261968 507134 262288 507218
rect 261968 506898 262010 507134
rect 262246 506898 262288 507134
rect 261968 506866 262288 506898
rect 292688 507454 293008 507486
rect 292688 507218 292730 507454
rect 292966 507218 293008 507454
rect 292688 507134 293008 507218
rect 292688 506898 292730 507134
rect 292966 506898 293008 507134
rect 292688 506866 293008 506898
rect 323408 507454 323728 507486
rect 323408 507218 323450 507454
rect 323686 507218 323728 507454
rect 323408 507134 323728 507218
rect 323408 506898 323450 507134
rect 323686 506898 323728 507134
rect 323408 506866 323728 506898
rect 354128 507454 354448 507486
rect 354128 507218 354170 507454
rect 354406 507218 354448 507454
rect 354128 507134 354448 507218
rect 354128 506898 354170 507134
rect 354406 506898 354448 507134
rect 354128 506866 354448 506898
rect 384848 507454 385168 507486
rect 384848 507218 384890 507454
rect 385126 507218 385168 507454
rect 384848 507134 385168 507218
rect 384848 506898 384890 507134
rect 385126 506898 385168 507134
rect 384848 506866 385168 506898
rect 415568 507454 415888 507486
rect 415568 507218 415610 507454
rect 415846 507218 415888 507454
rect 415568 507134 415888 507218
rect 415568 506898 415610 507134
rect 415846 506898 415888 507134
rect 415568 506866 415888 506898
rect 446288 507454 446608 507486
rect 446288 507218 446330 507454
rect 446566 507218 446608 507454
rect 446288 507134 446608 507218
rect 446288 506898 446330 507134
rect 446566 506898 446608 507134
rect 446288 506866 446608 506898
rect 477008 507454 477328 507486
rect 477008 507218 477050 507454
rect 477286 507218 477328 507454
rect 477008 507134 477328 507218
rect 477008 506898 477050 507134
rect 477286 506898 477328 507134
rect 477008 506866 477328 506898
rect 507728 507454 508048 507486
rect 507728 507218 507770 507454
rect 508006 507218 508048 507454
rect 507728 507134 508048 507218
rect 507728 506898 507770 507134
rect 508006 506898 508048 507134
rect 507728 506866 508048 506898
rect 538448 507454 538768 507486
rect 538448 507218 538490 507454
rect 538726 507218 538768 507454
rect 538448 507134 538768 507218
rect 538448 506898 538490 507134
rect 538726 506898 538768 507134
rect 538448 506866 538768 506898
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 31568 475174 31888 475206
rect 31568 474938 31610 475174
rect 31846 474938 31888 475174
rect 31568 474854 31888 474938
rect 31568 474618 31610 474854
rect 31846 474618 31888 474854
rect 31568 474586 31888 474618
rect 62288 475174 62608 475206
rect 62288 474938 62330 475174
rect 62566 474938 62608 475174
rect 62288 474854 62608 474938
rect 62288 474618 62330 474854
rect 62566 474618 62608 474854
rect 62288 474586 62608 474618
rect 93008 475174 93328 475206
rect 93008 474938 93050 475174
rect 93286 474938 93328 475174
rect 93008 474854 93328 474938
rect 93008 474618 93050 474854
rect 93286 474618 93328 474854
rect 93008 474586 93328 474618
rect 123728 475174 124048 475206
rect 123728 474938 123770 475174
rect 124006 474938 124048 475174
rect 123728 474854 124048 474938
rect 123728 474618 123770 474854
rect 124006 474618 124048 474854
rect 123728 474586 124048 474618
rect 154448 475174 154768 475206
rect 154448 474938 154490 475174
rect 154726 474938 154768 475174
rect 154448 474854 154768 474938
rect 154448 474618 154490 474854
rect 154726 474618 154768 474854
rect 154448 474586 154768 474618
rect 185168 475174 185488 475206
rect 185168 474938 185210 475174
rect 185446 474938 185488 475174
rect 185168 474854 185488 474938
rect 185168 474618 185210 474854
rect 185446 474618 185488 474854
rect 185168 474586 185488 474618
rect 215888 475174 216208 475206
rect 215888 474938 215930 475174
rect 216166 474938 216208 475174
rect 215888 474854 216208 474938
rect 215888 474618 215930 474854
rect 216166 474618 216208 474854
rect 215888 474586 216208 474618
rect 246608 475174 246928 475206
rect 246608 474938 246650 475174
rect 246886 474938 246928 475174
rect 246608 474854 246928 474938
rect 246608 474618 246650 474854
rect 246886 474618 246928 474854
rect 246608 474586 246928 474618
rect 277328 475174 277648 475206
rect 277328 474938 277370 475174
rect 277606 474938 277648 475174
rect 277328 474854 277648 474938
rect 277328 474618 277370 474854
rect 277606 474618 277648 474854
rect 277328 474586 277648 474618
rect 308048 475174 308368 475206
rect 308048 474938 308090 475174
rect 308326 474938 308368 475174
rect 308048 474854 308368 474938
rect 308048 474618 308090 474854
rect 308326 474618 308368 474854
rect 308048 474586 308368 474618
rect 338768 475174 339088 475206
rect 338768 474938 338810 475174
rect 339046 474938 339088 475174
rect 338768 474854 339088 474938
rect 338768 474618 338810 474854
rect 339046 474618 339088 474854
rect 338768 474586 339088 474618
rect 369488 475174 369808 475206
rect 369488 474938 369530 475174
rect 369766 474938 369808 475174
rect 369488 474854 369808 474938
rect 369488 474618 369530 474854
rect 369766 474618 369808 474854
rect 369488 474586 369808 474618
rect 400208 475174 400528 475206
rect 400208 474938 400250 475174
rect 400486 474938 400528 475174
rect 400208 474854 400528 474938
rect 400208 474618 400250 474854
rect 400486 474618 400528 474854
rect 400208 474586 400528 474618
rect 430928 475174 431248 475206
rect 430928 474938 430970 475174
rect 431206 474938 431248 475174
rect 430928 474854 431248 474938
rect 430928 474618 430970 474854
rect 431206 474618 431248 474854
rect 430928 474586 431248 474618
rect 461648 475174 461968 475206
rect 461648 474938 461690 475174
rect 461926 474938 461968 475174
rect 461648 474854 461968 474938
rect 461648 474618 461690 474854
rect 461926 474618 461968 474854
rect 461648 474586 461968 474618
rect 492368 475174 492688 475206
rect 492368 474938 492410 475174
rect 492646 474938 492688 475174
rect 492368 474854 492688 474938
rect 492368 474618 492410 474854
rect 492646 474618 492688 474854
rect 492368 474586 492688 474618
rect 523088 475174 523408 475206
rect 523088 474938 523130 475174
rect 523366 474938 523408 475174
rect 523088 474854 523408 474938
rect 523088 474618 523130 474854
rect 523366 474618 523408 474854
rect 523088 474586 523408 474618
rect 16208 471454 16528 471486
rect 16208 471218 16250 471454
rect 16486 471218 16528 471454
rect 16208 471134 16528 471218
rect 16208 470898 16250 471134
rect 16486 470898 16528 471134
rect 16208 470866 16528 470898
rect 46928 471454 47248 471486
rect 46928 471218 46970 471454
rect 47206 471218 47248 471454
rect 46928 471134 47248 471218
rect 46928 470898 46970 471134
rect 47206 470898 47248 471134
rect 46928 470866 47248 470898
rect 77648 471454 77968 471486
rect 77648 471218 77690 471454
rect 77926 471218 77968 471454
rect 77648 471134 77968 471218
rect 77648 470898 77690 471134
rect 77926 470898 77968 471134
rect 77648 470866 77968 470898
rect 108368 471454 108688 471486
rect 108368 471218 108410 471454
rect 108646 471218 108688 471454
rect 108368 471134 108688 471218
rect 108368 470898 108410 471134
rect 108646 470898 108688 471134
rect 108368 470866 108688 470898
rect 139088 471454 139408 471486
rect 139088 471218 139130 471454
rect 139366 471218 139408 471454
rect 139088 471134 139408 471218
rect 139088 470898 139130 471134
rect 139366 470898 139408 471134
rect 139088 470866 139408 470898
rect 169808 471454 170128 471486
rect 169808 471218 169850 471454
rect 170086 471218 170128 471454
rect 169808 471134 170128 471218
rect 169808 470898 169850 471134
rect 170086 470898 170128 471134
rect 169808 470866 170128 470898
rect 200528 471454 200848 471486
rect 200528 471218 200570 471454
rect 200806 471218 200848 471454
rect 200528 471134 200848 471218
rect 200528 470898 200570 471134
rect 200806 470898 200848 471134
rect 200528 470866 200848 470898
rect 231248 471454 231568 471486
rect 231248 471218 231290 471454
rect 231526 471218 231568 471454
rect 231248 471134 231568 471218
rect 231248 470898 231290 471134
rect 231526 470898 231568 471134
rect 231248 470866 231568 470898
rect 261968 471454 262288 471486
rect 261968 471218 262010 471454
rect 262246 471218 262288 471454
rect 261968 471134 262288 471218
rect 261968 470898 262010 471134
rect 262246 470898 262288 471134
rect 261968 470866 262288 470898
rect 292688 471454 293008 471486
rect 292688 471218 292730 471454
rect 292966 471218 293008 471454
rect 292688 471134 293008 471218
rect 292688 470898 292730 471134
rect 292966 470898 293008 471134
rect 292688 470866 293008 470898
rect 323408 471454 323728 471486
rect 323408 471218 323450 471454
rect 323686 471218 323728 471454
rect 323408 471134 323728 471218
rect 323408 470898 323450 471134
rect 323686 470898 323728 471134
rect 323408 470866 323728 470898
rect 354128 471454 354448 471486
rect 354128 471218 354170 471454
rect 354406 471218 354448 471454
rect 354128 471134 354448 471218
rect 354128 470898 354170 471134
rect 354406 470898 354448 471134
rect 354128 470866 354448 470898
rect 384848 471454 385168 471486
rect 384848 471218 384890 471454
rect 385126 471218 385168 471454
rect 384848 471134 385168 471218
rect 384848 470898 384890 471134
rect 385126 470898 385168 471134
rect 384848 470866 385168 470898
rect 415568 471454 415888 471486
rect 415568 471218 415610 471454
rect 415846 471218 415888 471454
rect 415568 471134 415888 471218
rect 415568 470898 415610 471134
rect 415846 470898 415888 471134
rect 415568 470866 415888 470898
rect 446288 471454 446608 471486
rect 446288 471218 446330 471454
rect 446566 471218 446608 471454
rect 446288 471134 446608 471218
rect 446288 470898 446330 471134
rect 446566 470898 446608 471134
rect 446288 470866 446608 470898
rect 477008 471454 477328 471486
rect 477008 471218 477050 471454
rect 477286 471218 477328 471454
rect 477008 471134 477328 471218
rect 477008 470898 477050 471134
rect 477286 470898 477328 471134
rect 477008 470866 477328 470898
rect 507728 471454 508048 471486
rect 507728 471218 507770 471454
rect 508006 471218 508048 471454
rect 507728 471134 508048 471218
rect 507728 470898 507770 471134
rect 508006 470898 508048 471134
rect 507728 470866 508048 470898
rect 538448 471454 538768 471486
rect 538448 471218 538490 471454
rect 538726 471218 538768 471454
rect 538448 471134 538768 471218
rect 538448 470898 538490 471134
rect 538726 470898 538768 471134
rect 538448 470866 538768 470898
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 31568 439174 31888 439206
rect 31568 438938 31610 439174
rect 31846 438938 31888 439174
rect 31568 438854 31888 438938
rect 31568 438618 31610 438854
rect 31846 438618 31888 438854
rect 31568 438586 31888 438618
rect 62288 439174 62608 439206
rect 62288 438938 62330 439174
rect 62566 438938 62608 439174
rect 62288 438854 62608 438938
rect 62288 438618 62330 438854
rect 62566 438618 62608 438854
rect 62288 438586 62608 438618
rect 93008 439174 93328 439206
rect 93008 438938 93050 439174
rect 93286 438938 93328 439174
rect 93008 438854 93328 438938
rect 93008 438618 93050 438854
rect 93286 438618 93328 438854
rect 93008 438586 93328 438618
rect 123728 439174 124048 439206
rect 123728 438938 123770 439174
rect 124006 438938 124048 439174
rect 123728 438854 124048 438938
rect 123728 438618 123770 438854
rect 124006 438618 124048 438854
rect 123728 438586 124048 438618
rect 154448 439174 154768 439206
rect 154448 438938 154490 439174
rect 154726 438938 154768 439174
rect 154448 438854 154768 438938
rect 154448 438618 154490 438854
rect 154726 438618 154768 438854
rect 154448 438586 154768 438618
rect 185168 439174 185488 439206
rect 185168 438938 185210 439174
rect 185446 438938 185488 439174
rect 185168 438854 185488 438938
rect 185168 438618 185210 438854
rect 185446 438618 185488 438854
rect 185168 438586 185488 438618
rect 215888 439174 216208 439206
rect 215888 438938 215930 439174
rect 216166 438938 216208 439174
rect 215888 438854 216208 438938
rect 215888 438618 215930 438854
rect 216166 438618 216208 438854
rect 215888 438586 216208 438618
rect 246608 439174 246928 439206
rect 246608 438938 246650 439174
rect 246886 438938 246928 439174
rect 246608 438854 246928 438938
rect 246608 438618 246650 438854
rect 246886 438618 246928 438854
rect 246608 438586 246928 438618
rect 277328 439174 277648 439206
rect 277328 438938 277370 439174
rect 277606 438938 277648 439174
rect 277328 438854 277648 438938
rect 277328 438618 277370 438854
rect 277606 438618 277648 438854
rect 277328 438586 277648 438618
rect 308048 439174 308368 439206
rect 308048 438938 308090 439174
rect 308326 438938 308368 439174
rect 308048 438854 308368 438938
rect 308048 438618 308090 438854
rect 308326 438618 308368 438854
rect 308048 438586 308368 438618
rect 338768 439174 339088 439206
rect 338768 438938 338810 439174
rect 339046 438938 339088 439174
rect 338768 438854 339088 438938
rect 338768 438618 338810 438854
rect 339046 438618 339088 438854
rect 338768 438586 339088 438618
rect 369488 439174 369808 439206
rect 369488 438938 369530 439174
rect 369766 438938 369808 439174
rect 369488 438854 369808 438938
rect 369488 438618 369530 438854
rect 369766 438618 369808 438854
rect 369488 438586 369808 438618
rect 400208 439174 400528 439206
rect 400208 438938 400250 439174
rect 400486 438938 400528 439174
rect 400208 438854 400528 438938
rect 400208 438618 400250 438854
rect 400486 438618 400528 438854
rect 400208 438586 400528 438618
rect 430928 439174 431248 439206
rect 430928 438938 430970 439174
rect 431206 438938 431248 439174
rect 430928 438854 431248 438938
rect 430928 438618 430970 438854
rect 431206 438618 431248 438854
rect 430928 438586 431248 438618
rect 461648 439174 461968 439206
rect 461648 438938 461690 439174
rect 461926 438938 461968 439174
rect 461648 438854 461968 438938
rect 461648 438618 461690 438854
rect 461926 438618 461968 438854
rect 461648 438586 461968 438618
rect 492368 439174 492688 439206
rect 492368 438938 492410 439174
rect 492646 438938 492688 439174
rect 492368 438854 492688 438938
rect 492368 438618 492410 438854
rect 492646 438618 492688 438854
rect 492368 438586 492688 438618
rect 523088 439174 523408 439206
rect 523088 438938 523130 439174
rect 523366 438938 523408 439174
rect 523088 438854 523408 438938
rect 523088 438618 523130 438854
rect 523366 438618 523408 438854
rect 523088 438586 523408 438618
rect 16208 435454 16528 435486
rect 16208 435218 16250 435454
rect 16486 435218 16528 435454
rect 16208 435134 16528 435218
rect 16208 434898 16250 435134
rect 16486 434898 16528 435134
rect 16208 434866 16528 434898
rect 46928 435454 47248 435486
rect 46928 435218 46970 435454
rect 47206 435218 47248 435454
rect 46928 435134 47248 435218
rect 46928 434898 46970 435134
rect 47206 434898 47248 435134
rect 46928 434866 47248 434898
rect 77648 435454 77968 435486
rect 77648 435218 77690 435454
rect 77926 435218 77968 435454
rect 77648 435134 77968 435218
rect 77648 434898 77690 435134
rect 77926 434898 77968 435134
rect 77648 434866 77968 434898
rect 108368 435454 108688 435486
rect 108368 435218 108410 435454
rect 108646 435218 108688 435454
rect 108368 435134 108688 435218
rect 108368 434898 108410 435134
rect 108646 434898 108688 435134
rect 108368 434866 108688 434898
rect 139088 435454 139408 435486
rect 139088 435218 139130 435454
rect 139366 435218 139408 435454
rect 139088 435134 139408 435218
rect 139088 434898 139130 435134
rect 139366 434898 139408 435134
rect 139088 434866 139408 434898
rect 169808 435454 170128 435486
rect 169808 435218 169850 435454
rect 170086 435218 170128 435454
rect 169808 435134 170128 435218
rect 169808 434898 169850 435134
rect 170086 434898 170128 435134
rect 169808 434866 170128 434898
rect 200528 435454 200848 435486
rect 200528 435218 200570 435454
rect 200806 435218 200848 435454
rect 200528 435134 200848 435218
rect 200528 434898 200570 435134
rect 200806 434898 200848 435134
rect 200528 434866 200848 434898
rect 231248 435454 231568 435486
rect 231248 435218 231290 435454
rect 231526 435218 231568 435454
rect 231248 435134 231568 435218
rect 231248 434898 231290 435134
rect 231526 434898 231568 435134
rect 231248 434866 231568 434898
rect 261968 435454 262288 435486
rect 261968 435218 262010 435454
rect 262246 435218 262288 435454
rect 261968 435134 262288 435218
rect 261968 434898 262010 435134
rect 262246 434898 262288 435134
rect 261968 434866 262288 434898
rect 292688 435454 293008 435486
rect 292688 435218 292730 435454
rect 292966 435218 293008 435454
rect 292688 435134 293008 435218
rect 292688 434898 292730 435134
rect 292966 434898 293008 435134
rect 292688 434866 293008 434898
rect 323408 435454 323728 435486
rect 323408 435218 323450 435454
rect 323686 435218 323728 435454
rect 323408 435134 323728 435218
rect 323408 434898 323450 435134
rect 323686 434898 323728 435134
rect 323408 434866 323728 434898
rect 354128 435454 354448 435486
rect 354128 435218 354170 435454
rect 354406 435218 354448 435454
rect 354128 435134 354448 435218
rect 354128 434898 354170 435134
rect 354406 434898 354448 435134
rect 354128 434866 354448 434898
rect 384848 435454 385168 435486
rect 384848 435218 384890 435454
rect 385126 435218 385168 435454
rect 384848 435134 385168 435218
rect 384848 434898 384890 435134
rect 385126 434898 385168 435134
rect 384848 434866 385168 434898
rect 415568 435454 415888 435486
rect 415568 435218 415610 435454
rect 415846 435218 415888 435454
rect 415568 435134 415888 435218
rect 415568 434898 415610 435134
rect 415846 434898 415888 435134
rect 415568 434866 415888 434898
rect 446288 435454 446608 435486
rect 446288 435218 446330 435454
rect 446566 435218 446608 435454
rect 446288 435134 446608 435218
rect 446288 434898 446330 435134
rect 446566 434898 446608 435134
rect 446288 434866 446608 434898
rect 477008 435454 477328 435486
rect 477008 435218 477050 435454
rect 477286 435218 477328 435454
rect 477008 435134 477328 435218
rect 477008 434898 477050 435134
rect 477286 434898 477328 435134
rect 477008 434866 477328 434898
rect 507728 435454 508048 435486
rect 507728 435218 507770 435454
rect 508006 435218 508048 435454
rect 507728 435134 508048 435218
rect 507728 434898 507770 435134
rect 508006 434898 508048 435134
rect 507728 434866 508048 434898
rect 538448 435454 538768 435486
rect 538448 435218 538490 435454
rect 538726 435218 538768 435454
rect 538448 435134 538768 435218
rect 538448 434898 538490 435134
rect 538726 434898 538768 435134
rect 538448 434866 538768 434898
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 31568 403174 31888 403206
rect 31568 402938 31610 403174
rect 31846 402938 31888 403174
rect 31568 402854 31888 402938
rect 31568 402618 31610 402854
rect 31846 402618 31888 402854
rect 31568 402586 31888 402618
rect 62288 403174 62608 403206
rect 62288 402938 62330 403174
rect 62566 402938 62608 403174
rect 62288 402854 62608 402938
rect 62288 402618 62330 402854
rect 62566 402618 62608 402854
rect 62288 402586 62608 402618
rect 93008 403174 93328 403206
rect 93008 402938 93050 403174
rect 93286 402938 93328 403174
rect 93008 402854 93328 402938
rect 93008 402618 93050 402854
rect 93286 402618 93328 402854
rect 93008 402586 93328 402618
rect 123728 403174 124048 403206
rect 123728 402938 123770 403174
rect 124006 402938 124048 403174
rect 123728 402854 124048 402938
rect 123728 402618 123770 402854
rect 124006 402618 124048 402854
rect 123728 402586 124048 402618
rect 154448 403174 154768 403206
rect 154448 402938 154490 403174
rect 154726 402938 154768 403174
rect 154448 402854 154768 402938
rect 154448 402618 154490 402854
rect 154726 402618 154768 402854
rect 154448 402586 154768 402618
rect 185168 403174 185488 403206
rect 185168 402938 185210 403174
rect 185446 402938 185488 403174
rect 185168 402854 185488 402938
rect 185168 402618 185210 402854
rect 185446 402618 185488 402854
rect 185168 402586 185488 402618
rect 215888 403174 216208 403206
rect 215888 402938 215930 403174
rect 216166 402938 216208 403174
rect 215888 402854 216208 402938
rect 215888 402618 215930 402854
rect 216166 402618 216208 402854
rect 215888 402586 216208 402618
rect 246608 403174 246928 403206
rect 246608 402938 246650 403174
rect 246886 402938 246928 403174
rect 246608 402854 246928 402938
rect 246608 402618 246650 402854
rect 246886 402618 246928 402854
rect 246608 402586 246928 402618
rect 277328 403174 277648 403206
rect 277328 402938 277370 403174
rect 277606 402938 277648 403174
rect 277328 402854 277648 402938
rect 277328 402618 277370 402854
rect 277606 402618 277648 402854
rect 277328 402586 277648 402618
rect 308048 403174 308368 403206
rect 308048 402938 308090 403174
rect 308326 402938 308368 403174
rect 308048 402854 308368 402938
rect 308048 402618 308090 402854
rect 308326 402618 308368 402854
rect 308048 402586 308368 402618
rect 338768 403174 339088 403206
rect 338768 402938 338810 403174
rect 339046 402938 339088 403174
rect 338768 402854 339088 402938
rect 338768 402618 338810 402854
rect 339046 402618 339088 402854
rect 338768 402586 339088 402618
rect 369488 403174 369808 403206
rect 369488 402938 369530 403174
rect 369766 402938 369808 403174
rect 369488 402854 369808 402938
rect 369488 402618 369530 402854
rect 369766 402618 369808 402854
rect 369488 402586 369808 402618
rect 400208 403174 400528 403206
rect 400208 402938 400250 403174
rect 400486 402938 400528 403174
rect 400208 402854 400528 402938
rect 400208 402618 400250 402854
rect 400486 402618 400528 402854
rect 400208 402586 400528 402618
rect 430928 403174 431248 403206
rect 430928 402938 430970 403174
rect 431206 402938 431248 403174
rect 430928 402854 431248 402938
rect 430928 402618 430970 402854
rect 431206 402618 431248 402854
rect 430928 402586 431248 402618
rect 461648 403174 461968 403206
rect 461648 402938 461690 403174
rect 461926 402938 461968 403174
rect 461648 402854 461968 402938
rect 461648 402618 461690 402854
rect 461926 402618 461968 402854
rect 461648 402586 461968 402618
rect 492368 403174 492688 403206
rect 492368 402938 492410 403174
rect 492646 402938 492688 403174
rect 492368 402854 492688 402938
rect 492368 402618 492410 402854
rect 492646 402618 492688 402854
rect 492368 402586 492688 402618
rect 523088 403174 523408 403206
rect 523088 402938 523130 403174
rect 523366 402938 523408 403174
rect 523088 402854 523408 402938
rect 523088 402618 523130 402854
rect 523366 402618 523408 402854
rect 523088 402586 523408 402618
rect 16208 399454 16528 399486
rect 16208 399218 16250 399454
rect 16486 399218 16528 399454
rect 16208 399134 16528 399218
rect 16208 398898 16250 399134
rect 16486 398898 16528 399134
rect 16208 398866 16528 398898
rect 46928 399454 47248 399486
rect 46928 399218 46970 399454
rect 47206 399218 47248 399454
rect 46928 399134 47248 399218
rect 46928 398898 46970 399134
rect 47206 398898 47248 399134
rect 46928 398866 47248 398898
rect 77648 399454 77968 399486
rect 77648 399218 77690 399454
rect 77926 399218 77968 399454
rect 77648 399134 77968 399218
rect 77648 398898 77690 399134
rect 77926 398898 77968 399134
rect 77648 398866 77968 398898
rect 108368 399454 108688 399486
rect 108368 399218 108410 399454
rect 108646 399218 108688 399454
rect 108368 399134 108688 399218
rect 108368 398898 108410 399134
rect 108646 398898 108688 399134
rect 108368 398866 108688 398898
rect 139088 399454 139408 399486
rect 139088 399218 139130 399454
rect 139366 399218 139408 399454
rect 139088 399134 139408 399218
rect 139088 398898 139130 399134
rect 139366 398898 139408 399134
rect 139088 398866 139408 398898
rect 169808 399454 170128 399486
rect 169808 399218 169850 399454
rect 170086 399218 170128 399454
rect 169808 399134 170128 399218
rect 169808 398898 169850 399134
rect 170086 398898 170128 399134
rect 169808 398866 170128 398898
rect 200528 399454 200848 399486
rect 200528 399218 200570 399454
rect 200806 399218 200848 399454
rect 200528 399134 200848 399218
rect 200528 398898 200570 399134
rect 200806 398898 200848 399134
rect 200528 398866 200848 398898
rect 231248 399454 231568 399486
rect 231248 399218 231290 399454
rect 231526 399218 231568 399454
rect 231248 399134 231568 399218
rect 231248 398898 231290 399134
rect 231526 398898 231568 399134
rect 231248 398866 231568 398898
rect 261968 399454 262288 399486
rect 261968 399218 262010 399454
rect 262246 399218 262288 399454
rect 261968 399134 262288 399218
rect 261968 398898 262010 399134
rect 262246 398898 262288 399134
rect 261968 398866 262288 398898
rect 292688 399454 293008 399486
rect 292688 399218 292730 399454
rect 292966 399218 293008 399454
rect 292688 399134 293008 399218
rect 292688 398898 292730 399134
rect 292966 398898 293008 399134
rect 292688 398866 293008 398898
rect 323408 399454 323728 399486
rect 323408 399218 323450 399454
rect 323686 399218 323728 399454
rect 323408 399134 323728 399218
rect 323408 398898 323450 399134
rect 323686 398898 323728 399134
rect 323408 398866 323728 398898
rect 354128 399454 354448 399486
rect 354128 399218 354170 399454
rect 354406 399218 354448 399454
rect 354128 399134 354448 399218
rect 354128 398898 354170 399134
rect 354406 398898 354448 399134
rect 354128 398866 354448 398898
rect 384848 399454 385168 399486
rect 384848 399218 384890 399454
rect 385126 399218 385168 399454
rect 384848 399134 385168 399218
rect 384848 398898 384890 399134
rect 385126 398898 385168 399134
rect 384848 398866 385168 398898
rect 415568 399454 415888 399486
rect 415568 399218 415610 399454
rect 415846 399218 415888 399454
rect 415568 399134 415888 399218
rect 415568 398898 415610 399134
rect 415846 398898 415888 399134
rect 415568 398866 415888 398898
rect 446288 399454 446608 399486
rect 446288 399218 446330 399454
rect 446566 399218 446608 399454
rect 446288 399134 446608 399218
rect 446288 398898 446330 399134
rect 446566 398898 446608 399134
rect 446288 398866 446608 398898
rect 477008 399454 477328 399486
rect 477008 399218 477050 399454
rect 477286 399218 477328 399454
rect 477008 399134 477328 399218
rect 477008 398898 477050 399134
rect 477286 398898 477328 399134
rect 477008 398866 477328 398898
rect 507728 399454 508048 399486
rect 507728 399218 507770 399454
rect 508006 399218 508048 399454
rect 507728 399134 508048 399218
rect 507728 398898 507770 399134
rect 508006 398898 508048 399134
rect 507728 398866 508048 398898
rect 538448 399454 538768 399486
rect 538448 399218 538490 399454
rect 538726 399218 538768 399454
rect 538448 399134 538768 399218
rect 538448 398898 538490 399134
rect 538726 398898 538768 399134
rect 538448 398866 538768 398898
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 556674 378334 557294 413778
rect 556674 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 557294 378334
rect 556674 378014 557294 378098
rect 556674 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 557294 378014
rect 31568 367174 31888 367206
rect 31568 366938 31610 367174
rect 31846 366938 31888 367174
rect 31568 366854 31888 366938
rect 31568 366618 31610 366854
rect 31846 366618 31888 366854
rect 31568 366586 31888 366618
rect 62288 367174 62608 367206
rect 62288 366938 62330 367174
rect 62566 366938 62608 367174
rect 62288 366854 62608 366938
rect 62288 366618 62330 366854
rect 62566 366618 62608 366854
rect 62288 366586 62608 366618
rect 93008 367174 93328 367206
rect 93008 366938 93050 367174
rect 93286 366938 93328 367174
rect 93008 366854 93328 366938
rect 93008 366618 93050 366854
rect 93286 366618 93328 366854
rect 93008 366586 93328 366618
rect 123728 367174 124048 367206
rect 123728 366938 123770 367174
rect 124006 366938 124048 367174
rect 123728 366854 124048 366938
rect 123728 366618 123770 366854
rect 124006 366618 124048 366854
rect 123728 366586 124048 366618
rect 154448 367174 154768 367206
rect 154448 366938 154490 367174
rect 154726 366938 154768 367174
rect 154448 366854 154768 366938
rect 154448 366618 154490 366854
rect 154726 366618 154768 366854
rect 154448 366586 154768 366618
rect 185168 367174 185488 367206
rect 185168 366938 185210 367174
rect 185446 366938 185488 367174
rect 185168 366854 185488 366938
rect 185168 366618 185210 366854
rect 185446 366618 185488 366854
rect 185168 366586 185488 366618
rect 215888 367174 216208 367206
rect 215888 366938 215930 367174
rect 216166 366938 216208 367174
rect 215888 366854 216208 366938
rect 215888 366618 215930 366854
rect 216166 366618 216208 366854
rect 215888 366586 216208 366618
rect 246608 367174 246928 367206
rect 246608 366938 246650 367174
rect 246886 366938 246928 367174
rect 246608 366854 246928 366938
rect 246608 366618 246650 366854
rect 246886 366618 246928 366854
rect 246608 366586 246928 366618
rect 277328 367174 277648 367206
rect 277328 366938 277370 367174
rect 277606 366938 277648 367174
rect 277328 366854 277648 366938
rect 277328 366618 277370 366854
rect 277606 366618 277648 366854
rect 277328 366586 277648 366618
rect 308048 367174 308368 367206
rect 308048 366938 308090 367174
rect 308326 366938 308368 367174
rect 308048 366854 308368 366938
rect 308048 366618 308090 366854
rect 308326 366618 308368 366854
rect 308048 366586 308368 366618
rect 338768 367174 339088 367206
rect 338768 366938 338810 367174
rect 339046 366938 339088 367174
rect 338768 366854 339088 366938
rect 338768 366618 338810 366854
rect 339046 366618 339088 366854
rect 338768 366586 339088 366618
rect 369488 367174 369808 367206
rect 369488 366938 369530 367174
rect 369766 366938 369808 367174
rect 369488 366854 369808 366938
rect 369488 366618 369530 366854
rect 369766 366618 369808 366854
rect 369488 366586 369808 366618
rect 400208 367174 400528 367206
rect 400208 366938 400250 367174
rect 400486 366938 400528 367174
rect 400208 366854 400528 366938
rect 400208 366618 400250 366854
rect 400486 366618 400528 366854
rect 400208 366586 400528 366618
rect 430928 367174 431248 367206
rect 430928 366938 430970 367174
rect 431206 366938 431248 367174
rect 430928 366854 431248 366938
rect 430928 366618 430970 366854
rect 431206 366618 431248 366854
rect 430928 366586 431248 366618
rect 461648 367174 461968 367206
rect 461648 366938 461690 367174
rect 461926 366938 461968 367174
rect 461648 366854 461968 366938
rect 461648 366618 461690 366854
rect 461926 366618 461968 366854
rect 461648 366586 461968 366618
rect 492368 367174 492688 367206
rect 492368 366938 492410 367174
rect 492646 366938 492688 367174
rect 492368 366854 492688 366938
rect 492368 366618 492410 366854
rect 492646 366618 492688 366854
rect 492368 366586 492688 366618
rect 523088 367174 523408 367206
rect 523088 366938 523130 367174
rect 523366 366938 523408 367174
rect 523088 366854 523408 366938
rect 523088 366618 523130 366854
rect 523366 366618 523408 366854
rect 523088 366586 523408 366618
rect 16208 363454 16528 363486
rect 16208 363218 16250 363454
rect 16486 363218 16528 363454
rect 16208 363134 16528 363218
rect 16208 362898 16250 363134
rect 16486 362898 16528 363134
rect 16208 362866 16528 362898
rect 46928 363454 47248 363486
rect 46928 363218 46970 363454
rect 47206 363218 47248 363454
rect 46928 363134 47248 363218
rect 46928 362898 46970 363134
rect 47206 362898 47248 363134
rect 46928 362866 47248 362898
rect 77648 363454 77968 363486
rect 77648 363218 77690 363454
rect 77926 363218 77968 363454
rect 77648 363134 77968 363218
rect 77648 362898 77690 363134
rect 77926 362898 77968 363134
rect 77648 362866 77968 362898
rect 108368 363454 108688 363486
rect 108368 363218 108410 363454
rect 108646 363218 108688 363454
rect 108368 363134 108688 363218
rect 108368 362898 108410 363134
rect 108646 362898 108688 363134
rect 108368 362866 108688 362898
rect 139088 363454 139408 363486
rect 139088 363218 139130 363454
rect 139366 363218 139408 363454
rect 139088 363134 139408 363218
rect 139088 362898 139130 363134
rect 139366 362898 139408 363134
rect 139088 362866 139408 362898
rect 169808 363454 170128 363486
rect 169808 363218 169850 363454
rect 170086 363218 170128 363454
rect 169808 363134 170128 363218
rect 169808 362898 169850 363134
rect 170086 362898 170128 363134
rect 169808 362866 170128 362898
rect 200528 363454 200848 363486
rect 200528 363218 200570 363454
rect 200806 363218 200848 363454
rect 200528 363134 200848 363218
rect 200528 362898 200570 363134
rect 200806 362898 200848 363134
rect 200528 362866 200848 362898
rect 231248 363454 231568 363486
rect 231248 363218 231290 363454
rect 231526 363218 231568 363454
rect 231248 363134 231568 363218
rect 231248 362898 231290 363134
rect 231526 362898 231568 363134
rect 231248 362866 231568 362898
rect 261968 363454 262288 363486
rect 261968 363218 262010 363454
rect 262246 363218 262288 363454
rect 261968 363134 262288 363218
rect 261968 362898 262010 363134
rect 262246 362898 262288 363134
rect 261968 362866 262288 362898
rect 292688 363454 293008 363486
rect 292688 363218 292730 363454
rect 292966 363218 293008 363454
rect 292688 363134 293008 363218
rect 292688 362898 292730 363134
rect 292966 362898 293008 363134
rect 292688 362866 293008 362898
rect 323408 363454 323728 363486
rect 323408 363218 323450 363454
rect 323686 363218 323728 363454
rect 323408 363134 323728 363218
rect 323408 362898 323450 363134
rect 323686 362898 323728 363134
rect 323408 362866 323728 362898
rect 354128 363454 354448 363486
rect 354128 363218 354170 363454
rect 354406 363218 354448 363454
rect 354128 363134 354448 363218
rect 354128 362898 354170 363134
rect 354406 362898 354448 363134
rect 354128 362866 354448 362898
rect 384848 363454 385168 363486
rect 384848 363218 384890 363454
rect 385126 363218 385168 363454
rect 384848 363134 385168 363218
rect 384848 362898 384890 363134
rect 385126 362898 385168 363134
rect 384848 362866 385168 362898
rect 415568 363454 415888 363486
rect 415568 363218 415610 363454
rect 415846 363218 415888 363454
rect 415568 363134 415888 363218
rect 415568 362898 415610 363134
rect 415846 362898 415888 363134
rect 415568 362866 415888 362898
rect 446288 363454 446608 363486
rect 446288 363218 446330 363454
rect 446566 363218 446608 363454
rect 446288 363134 446608 363218
rect 446288 362898 446330 363134
rect 446566 362898 446608 363134
rect 446288 362866 446608 362898
rect 477008 363454 477328 363486
rect 477008 363218 477050 363454
rect 477286 363218 477328 363454
rect 477008 363134 477328 363218
rect 477008 362898 477050 363134
rect 477286 362898 477328 363134
rect 477008 362866 477328 362898
rect 507728 363454 508048 363486
rect 507728 363218 507770 363454
rect 508006 363218 508048 363454
rect 507728 363134 508048 363218
rect 507728 362898 507770 363134
rect 508006 362898 508048 363134
rect 507728 362866 508048 362898
rect 538448 363454 538768 363486
rect 538448 363218 538490 363454
rect 538726 363218 538768 363454
rect 538448 363134 538768 363218
rect 538448 362898 538490 363134
rect 538726 362898 538768 363134
rect 538448 362866 538768 362898
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 556674 342334 557294 377778
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 31568 331174 31888 331206
rect 31568 330938 31610 331174
rect 31846 330938 31888 331174
rect 31568 330854 31888 330938
rect 31568 330618 31610 330854
rect 31846 330618 31888 330854
rect 31568 330586 31888 330618
rect 62288 331174 62608 331206
rect 62288 330938 62330 331174
rect 62566 330938 62608 331174
rect 62288 330854 62608 330938
rect 62288 330618 62330 330854
rect 62566 330618 62608 330854
rect 62288 330586 62608 330618
rect 93008 331174 93328 331206
rect 93008 330938 93050 331174
rect 93286 330938 93328 331174
rect 93008 330854 93328 330938
rect 93008 330618 93050 330854
rect 93286 330618 93328 330854
rect 93008 330586 93328 330618
rect 123728 331174 124048 331206
rect 123728 330938 123770 331174
rect 124006 330938 124048 331174
rect 123728 330854 124048 330938
rect 123728 330618 123770 330854
rect 124006 330618 124048 330854
rect 123728 330586 124048 330618
rect 154448 331174 154768 331206
rect 154448 330938 154490 331174
rect 154726 330938 154768 331174
rect 154448 330854 154768 330938
rect 154448 330618 154490 330854
rect 154726 330618 154768 330854
rect 154448 330586 154768 330618
rect 185168 331174 185488 331206
rect 185168 330938 185210 331174
rect 185446 330938 185488 331174
rect 185168 330854 185488 330938
rect 185168 330618 185210 330854
rect 185446 330618 185488 330854
rect 185168 330586 185488 330618
rect 215888 331174 216208 331206
rect 215888 330938 215930 331174
rect 216166 330938 216208 331174
rect 215888 330854 216208 330938
rect 215888 330618 215930 330854
rect 216166 330618 216208 330854
rect 215888 330586 216208 330618
rect 246608 331174 246928 331206
rect 246608 330938 246650 331174
rect 246886 330938 246928 331174
rect 246608 330854 246928 330938
rect 246608 330618 246650 330854
rect 246886 330618 246928 330854
rect 246608 330586 246928 330618
rect 277328 331174 277648 331206
rect 277328 330938 277370 331174
rect 277606 330938 277648 331174
rect 277328 330854 277648 330938
rect 277328 330618 277370 330854
rect 277606 330618 277648 330854
rect 277328 330586 277648 330618
rect 308048 331174 308368 331206
rect 308048 330938 308090 331174
rect 308326 330938 308368 331174
rect 308048 330854 308368 330938
rect 308048 330618 308090 330854
rect 308326 330618 308368 330854
rect 308048 330586 308368 330618
rect 338768 331174 339088 331206
rect 338768 330938 338810 331174
rect 339046 330938 339088 331174
rect 338768 330854 339088 330938
rect 338768 330618 338810 330854
rect 339046 330618 339088 330854
rect 338768 330586 339088 330618
rect 369488 331174 369808 331206
rect 369488 330938 369530 331174
rect 369766 330938 369808 331174
rect 369488 330854 369808 330938
rect 369488 330618 369530 330854
rect 369766 330618 369808 330854
rect 369488 330586 369808 330618
rect 400208 331174 400528 331206
rect 400208 330938 400250 331174
rect 400486 330938 400528 331174
rect 400208 330854 400528 330938
rect 400208 330618 400250 330854
rect 400486 330618 400528 330854
rect 400208 330586 400528 330618
rect 430928 331174 431248 331206
rect 430928 330938 430970 331174
rect 431206 330938 431248 331174
rect 430928 330854 431248 330938
rect 430928 330618 430970 330854
rect 431206 330618 431248 330854
rect 430928 330586 431248 330618
rect 461648 331174 461968 331206
rect 461648 330938 461690 331174
rect 461926 330938 461968 331174
rect 461648 330854 461968 330938
rect 461648 330618 461690 330854
rect 461926 330618 461968 330854
rect 461648 330586 461968 330618
rect 492368 331174 492688 331206
rect 492368 330938 492410 331174
rect 492646 330938 492688 331174
rect 492368 330854 492688 330938
rect 492368 330618 492410 330854
rect 492646 330618 492688 330854
rect 492368 330586 492688 330618
rect 523088 331174 523408 331206
rect 523088 330938 523130 331174
rect 523366 330938 523408 331174
rect 523088 330854 523408 330938
rect 523088 330618 523130 330854
rect 523366 330618 523408 330854
rect 523088 330586 523408 330618
rect 16208 327454 16528 327486
rect 16208 327218 16250 327454
rect 16486 327218 16528 327454
rect 16208 327134 16528 327218
rect 16208 326898 16250 327134
rect 16486 326898 16528 327134
rect 16208 326866 16528 326898
rect 46928 327454 47248 327486
rect 46928 327218 46970 327454
rect 47206 327218 47248 327454
rect 46928 327134 47248 327218
rect 46928 326898 46970 327134
rect 47206 326898 47248 327134
rect 46928 326866 47248 326898
rect 77648 327454 77968 327486
rect 77648 327218 77690 327454
rect 77926 327218 77968 327454
rect 77648 327134 77968 327218
rect 77648 326898 77690 327134
rect 77926 326898 77968 327134
rect 77648 326866 77968 326898
rect 108368 327454 108688 327486
rect 108368 327218 108410 327454
rect 108646 327218 108688 327454
rect 108368 327134 108688 327218
rect 108368 326898 108410 327134
rect 108646 326898 108688 327134
rect 108368 326866 108688 326898
rect 139088 327454 139408 327486
rect 139088 327218 139130 327454
rect 139366 327218 139408 327454
rect 139088 327134 139408 327218
rect 139088 326898 139130 327134
rect 139366 326898 139408 327134
rect 139088 326866 139408 326898
rect 169808 327454 170128 327486
rect 169808 327218 169850 327454
rect 170086 327218 170128 327454
rect 169808 327134 170128 327218
rect 169808 326898 169850 327134
rect 170086 326898 170128 327134
rect 169808 326866 170128 326898
rect 200528 327454 200848 327486
rect 200528 327218 200570 327454
rect 200806 327218 200848 327454
rect 200528 327134 200848 327218
rect 200528 326898 200570 327134
rect 200806 326898 200848 327134
rect 200528 326866 200848 326898
rect 231248 327454 231568 327486
rect 231248 327218 231290 327454
rect 231526 327218 231568 327454
rect 231248 327134 231568 327218
rect 231248 326898 231290 327134
rect 231526 326898 231568 327134
rect 231248 326866 231568 326898
rect 261968 327454 262288 327486
rect 261968 327218 262010 327454
rect 262246 327218 262288 327454
rect 261968 327134 262288 327218
rect 261968 326898 262010 327134
rect 262246 326898 262288 327134
rect 261968 326866 262288 326898
rect 292688 327454 293008 327486
rect 292688 327218 292730 327454
rect 292966 327218 293008 327454
rect 292688 327134 293008 327218
rect 292688 326898 292730 327134
rect 292966 326898 293008 327134
rect 292688 326866 293008 326898
rect 323408 327454 323728 327486
rect 323408 327218 323450 327454
rect 323686 327218 323728 327454
rect 323408 327134 323728 327218
rect 323408 326898 323450 327134
rect 323686 326898 323728 327134
rect 323408 326866 323728 326898
rect 354128 327454 354448 327486
rect 354128 327218 354170 327454
rect 354406 327218 354448 327454
rect 354128 327134 354448 327218
rect 354128 326898 354170 327134
rect 354406 326898 354448 327134
rect 354128 326866 354448 326898
rect 384848 327454 385168 327486
rect 384848 327218 384890 327454
rect 385126 327218 385168 327454
rect 384848 327134 385168 327218
rect 384848 326898 384890 327134
rect 385126 326898 385168 327134
rect 384848 326866 385168 326898
rect 415568 327454 415888 327486
rect 415568 327218 415610 327454
rect 415846 327218 415888 327454
rect 415568 327134 415888 327218
rect 415568 326898 415610 327134
rect 415846 326898 415888 327134
rect 415568 326866 415888 326898
rect 446288 327454 446608 327486
rect 446288 327218 446330 327454
rect 446566 327218 446608 327454
rect 446288 327134 446608 327218
rect 446288 326898 446330 327134
rect 446566 326898 446608 327134
rect 446288 326866 446608 326898
rect 477008 327454 477328 327486
rect 477008 327218 477050 327454
rect 477286 327218 477328 327454
rect 477008 327134 477328 327218
rect 477008 326898 477050 327134
rect 477286 326898 477328 327134
rect 477008 326866 477328 326898
rect 507728 327454 508048 327486
rect 507728 327218 507770 327454
rect 508006 327218 508048 327454
rect 507728 327134 508048 327218
rect 507728 326898 507770 327134
rect 508006 326898 508048 327134
rect 507728 326866 508048 326898
rect 538448 327454 538768 327486
rect 538448 327218 538490 327454
rect 538726 327218 538768 327454
rect 538448 327134 538768 327218
rect 538448 326898 538490 327134
rect 538726 326898 538768 327134
rect 538448 326866 538768 326898
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 556674 306334 557294 341778
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 31568 295174 31888 295206
rect 31568 294938 31610 295174
rect 31846 294938 31888 295174
rect 31568 294854 31888 294938
rect 31568 294618 31610 294854
rect 31846 294618 31888 294854
rect 31568 294586 31888 294618
rect 62288 295174 62608 295206
rect 62288 294938 62330 295174
rect 62566 294938 62608 295174
rect 62288 294854 62608 294938
rect 62288 294618 62330 294854
rect 62566 294618 62608 294854
rect 62288 294586 62608 294618
rect 93008 295174 93328 295206
rect 93008 294938 93050 295174
rect 93286 294938 93328 295174
rect 93008 294854 93328 294938
rect 93008 294618 93050 294854
rect 93286 294618 93328 294854
rect 93008 294586 93328 294618
rect 123728 295174 124048 295206
rect 123728 294938 123770 295174
rect 124006 294938 124048 295174
rect 123728 294854 124048 294938
rect 123728 294618 123770 294854
rect 124006 294618 124048 294854
rect 123728 294586 124048 294618
rect 154448 295174 154768 295206
rect 154448 294938 154490 295174
rect 154726 294938 154768 295174
rect 154448 294854 154768 294938
rect 154448 294618 154490 294854
rect 154726 294618 154768 294854
rect 154448 294586 154768 294618
rect 185168 295174 185488 295206
rect 185168 294938 185210 295174
rect 185446 294938 185488 295174
rect 185168 294854 185488 294938
rect 185168 294618 185210 294854
rect 185446 294618 185488 294854
rect 185168 294586 185488 294618
rect 215888 295174 216208 295206
rect 215888 294938 215930 295174
rect 216166 294938 216208 295174
rect 215888 294854 216208 294938
rect 215888 294618 215930 294854
rect 216166 294618 216208 294854
rect 215888 294586 216208 294618
rect 246608 295174 246928 295206
rect 246608 294938 246650 295174
rect 246886 294938 246928 295174
rect 246608 294854 246928 294938
rect 246608 294618 246650 294854
rect 246886 294618 246928 294854
rect 246608 294586 246928 294618
rect 277328 295174 277648 295206
rect 277328 294938 277370 295174
rect 277606 294938 277648 295174
rect 277328 294854 277648 294938
rect 277328 294618 277370 294854
rect 277606 294618 277648 294854
rect 277328 294586 277648 294618
rect 308048 295174 308368 295206
rect 308048 294938 308090 295174
rect 308326 294938 308368 295174
rect 308048 294854 308368 294938
rect 308048 294618 308090 294854
rect 308326 294618 308368 294854
rect 308048 294586 308368 294618
rect 338768 295174 339088 295206
rect 338768 294938 338810 295174
rect 339046 294938 339088 295174
rect 338768 294854 339088 294938
rect 338768 294618 338810 294854
rect 339046 294618 339088 294854
rect 338768 294586 339088 294618
rect 369488 295174 369808 295206
rect 369488 294938 369530 295174
rect 369766 294938 369808 295174
rect 369488 294854 369808 294938
rect 369488 294618 369530 294854
rect 369766 294618 369808 294854
rect 369488 294586 369808 294618
rect 400208 295174 400528 295206
rect 400208 294938 400250 295174
rect 400486 294938 400528 295174
rect 400208 294854 400528 294938
rect 400208 294618 400250 294854
rect 400486 294618 400528 294854
rect 400208 294586 400528 294618
rect 430928 295174 431248 295206
rect 430928 294938 430970 295174
rect 431206 294938 431248 295174
rect 430928 294854 431248 294938
rect 430928 294618 430970 294854
rect 431206 294618 431248 294854
rect 430928 294586 431248 294618
rect 461648 295174 461968 295206
rect 461648 294938 461690 295174
rect 461926 294938 461968 295174
rect 461648 294854 461968 294938
rect 461648 294618 461690 294854
rect 461926 294618 461968 294854
rect 461648 294586 461968 294618
rect 492368 295174 492688 295206
rect 492368 294938 492410 295174
rect 492646 294938 492688 295174
rect 492368 294854 492688 294938
rect 492368 294618 492410 294854
rect 492646 294618 492688 294854
rect 492368 294586 492688 294618
rect 523088 295174 523408 295206
rect 523088 294938 523130 295174
rect 523366 294938 523408 295174
rect 523088 294854 523408 294938
rect 523088 294618 523130 294854
rect 523366 294618 523408 294854
rect 523088 294586 523408 294618
rect 16208 291454 16528 291486
rect 16208 291218 16250 291454
rect 16486 291218 16528 291454
rect 16208 291134 16528 291218
rect 16208 290898 16250 291134
rect 16486 290898 16528 291134
rect 16208 290866 16528 290898
rect 46928 291454 47248 291486
rect 46928 291218 46970 291454
rect 47206 291218 47248 291454
rect 46928 291134 47248 291218
rect 46928 290898 46970 291134
rect 47206 290898 47248 291134
rect 46928 290866 47248 290898
rect 77648 291454 77968 291486
rect 77648 291218 77690 291454
rect 77926 291218 77968 291454
rect 77648 291134 77968 291218
rect 77648 290898 77690 291134
rect 77926 290898 77968 291134
rect 77648 290866 77968 290898
rect 108368 291454 108688 291486
rect 108368 291218 108410 291454
rect 108646 291218 108688 291454
rect 108368 291134 108688 291218
rect 108368 290898 108410 291134
rect 108646 290898 108688 291134
rect 108368 290866 108688 290898
rect 139088 291454 139408 291486
rect 139088 291218 139130 291454
rect 139366 291218 139408 291454
rect 139088 291134 139408 291218
rect 139088 290898 139130 291134
rect 139366 290898 139408 291134
rect 139088 290866 139408 290898
rect 169808 291454 170128 291486
rect 169808 291218 169850 291454
rect 170086 291218 170128 291454
rect 169808 291134 170128 291218
rect 169808 290898 169850 291134
rect 170086 290898 170128 291134
rect 169808 290866 170128 290898
rect 200528 291454 200848 291486
rect 200528 291218 200570 291454
rect 200806 291218 200848 291454
rect 200528 291134 200848 291218
rect 200528 290898 200570 291134
rect 200806 290898 200848 291134
rect 200528 290866 200848 290898
rect 231248 291454 231568 291486
rect 231248 291218 231290 291454
rect 231526 291218 231568 291454
rect 231248 291134 231568 291218
rect 231248 290898 231290 291134
rect 231526 290898 231568 291134
rect 231248 290866 231568 290898
rect 261968 291454 262288 291486
rect 261968 291218 262010 291454
rect 262246 291218 262288 291454
rect 261968 291134 262288 291218
rect 261968 290898 262010 291134
rect 262246 290898 262288 291134
rect 261968 290866 262288 290898
rect 292688 291454 293008 291486
rect 292688 291218 292730 291454
rect 292966 291218 293008 291454
rect 292688 291134 293008 291218
rect 292688 290898 292730 291134
rect 292966 290898 293008 291134
rect 292688 290866 293008 290898
rect 323408 291454 323728 291486
rect 323408 291218 323450 291454
rect 323686 291218 323728 291454
rect 323408 291134 323728 291218
rect 323408 290898 323450 291134
rect 323686 290898 323728 291134
rect 323408 290866 323728 290898
rect 354128 291454 354448 291486
rect 354128 291218 354170 291454
rect 354406 291218 354448 291454
rect 354128 291134 354448 291218
rect 354128 290898 354170 291134
rect 354406 290898 354448 291134
rect 354128 290866 354448 290898
rect 384848 291454 385168 291486
rect 384848 291218 384890 291454
rect 385126 291218 385168 291454
rect 384848 291134 385168 291218
rect 384848 290898 384890 291134
rect 385126 290898 385168 291134
rect 384848 290866 385168 290898
rect 415568 291454 415888 291486
rect 415568 291218 415610 291454
rect 415846 291218 415888 291454
rect 415568 291134 415888 291218
rect 415568 290898 415610 291134
rect 415846 290898 415888 291134
rect 415568 290866 415888 290898
rect 446288 291454 446608 291486
rect 446288 291218 446330 291454
rect 446566 291218 446608 291454
rect 446288 291134 446608 291218
rect 446288 290898 446330 291134
rect 446566 290898 446608 291134
rect 446288 290866 446608 290898
rect 477008 291454 477328 291486
rect 477008 291218 477050 291454
rect 477286 291218 477328 291454
rect 477008 291134 477328 291218
rect 477008 290898 477050 291134
rect 477286 290898 477328 291134
rect 477008 290866 477328 290898
rect 507728 291454 508048 291486
rect 507728 291218 507770 291454
rect 508006 291218 508048 291454
rect 507728 291134 508048 291218
rect 507728 290898 507770 291134
rect 508006 290898 508048 291134
rect 507728 290866 508048 290898
rect 538448 291454 538768 291486
rect 538448 291218 538490 291454
rect 538726 291218 538768 291454
rect 538448 291134 538768 291218
rect 538448 290898 538490 291134
rect 538726 290898 538768 291134
rect 538448 290866 538768 290898
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 31568 259174 31888 259206
rect 31568 258938 31610 259174
rect 31846 258938 31888 259174
rect 31568 258854 31888 258938
rect 31568 258618 31610 258854
rect 31846 258618 31888 258854
rect 31568 258586 31888 258618
rect 62288 259174 62608 259206
rect 62288 258938 62330 259174
rect 62566 258938 62608 259174
rect 62288 258854 62608 258938
rect 62288 258618 62330 258854
rect 62566 258618 62608 258854
rect 62288 258586 62608 258618
rect 93008 259174 93328 259206
rect 93008 258938 93050 259174
rect 93286 258938 93328 259174
rect 93008 258854 93328 258938
rect 93008 258618 93050 258854
rect 93286 258618 93328 258854
rect 93008 258586 93328 258618
rect 123728 259174 124048 259206
rect 123728 258938 123770 259174
rect 124006 258938 124048 259174
rect 123728 258854 124048 258938
rect 123728 258618 123770 258854
rect 124006 258618 124048 258854
rect 123728 258586 124048 258618
rect 154448 259174 154768 259206
rect 154448 258938 154490 259174
rect 154726 258938 154768 259174
rect 154448 258854 154768 258938
rect 154448 258618 154490 258854
rect 154726 258618 154768 258854
rect 154448 258586 154768 258618
rect 185168 259174 185488 259206
rect 185168 258938 185210 259174
rect 185446 258938 185488 259174
rect 185168 258854 185488 258938
rect 185168 258618 185210 258854
rect 185446 258618 185488 258854
rect 185168 258586 185488 258618
rect 215888 259174 216208 259206
rect 215888 258938 215930 259174
rect 216166 258938 216208 259174
rect 215888 258854 216208 258938
rect 215888 258618 215930 258854
rect 216166 258618 216208 258854
rect 215888 258586 216208 258618
rect 246608 259174 246928 259206
rect 246608 258938 246650 259174
rect 246886 258938 246928 259174
rect 246608 258854 246928 258938
rect 246608 258618 246650 258854
rect 246886 258618 246928 258854
rect 246608 258586 246928 258618
rect 277328 259174 277648 259206
rect 277328 258938 277370 259174
rect 277606 258938 277648 259174
rect 277328 258854 277648 258938
rect 277328 258618 277370 258854
rect 277606 258618 277648 258854
rect 277328 258586 277648 258618
rect 308048 259174 308368 259206
rect 308048 258938 308090 259174
rect 308326 258938 308368 259174
rect 308048 258854 308368 258938
rect 308048 258618 308090 258854
rect 308326 258618 308368 258854
rect 308048 258586 308368 258618
rect 338768 259174 339088 259206
rect 338768 258938 338810 259174
rect 339046 258938 339088 259174
rect 338768 258854 339088 258938
rect 338768 258618 338810 258854
rect 339046 258618 339088 258854
rect 338768 258586 339088 258618
rect 369488 259174 369808 259206
rect 369488 258938 369530 259174
rect 369766 258938 369808 259174
rect 369488 258854 369808 258938
rect 369488 258618 369530 258854
rect 369766 258618 369808 258854
rect 369488 258586 369808 258618
rect 400208 259174 400528 259206
rect 400208 258938 400250 259174
rect 400486 258938 400528 259174
rect 400208 258854 400528 258938
rect 400208 258618 400250 258854
rect 400486 258618 400528 258854
rect 400208 258586 400528 258618
rect 430928 259174 431248 259206
rect 430928 258938 430970 259174
rect 431206 258938 431248 259174
rect 430928 258854 431248 258938
rect 430928 258618 430970 258854
rect 431206 258618 431248 258854
rect 430928 258586 431248 258618
rect 461648 259174 461968 259206
rect 461648 258938 461690 259174
rect 461926 258938 461968 259174
rect 461648 258854 461968 258938
rect 461648 258618 461690 258854
rect 461926 258618 461968 258854
rect 461648 258586 461968 258618
rect 492368 259174 492688 259206
rect 492368 258938 492410 259174
rect 492646 258938 492688 259174
rect 492368 258854 492688 258938
rect 492368 258618 492410 258854
rect 492646 258618 492688 258854
rect 492368 258586 492688 258618
rect 523088 259174 523408 259206
rect 523088 258938 523130 259174
rect 523366 258938 523408 259174
rect 523088 258854 523408 258938
rect 523088 258618 523130 258854
rect 523366 258618 523408 258854
rect 523088 258586 523408 258618
rect 16208 255454 16528 255486
rect 16208 255218 16250 255454
rect 16486 255218 16528 255454
rect 16208 255134 16528 255218
rect 16208 254898 16250 255134
rect 16486 254898 16528 255134
rect 16208 254866 16528 254898
rect 46928 255454 47248 255486
rect 46928 255218 46970 255454
rect 47206 255218 47248 255454
rect 46928 255134 47248 255218
rect 46928 254898 46970 255134
rect 47206 254898 47248 255134
rect 46928 254866 47248 254898
rect 77648 255454 77968 255486
rect 77648 255218 77690 255454
rect 77926 255218 77968 255454
rect 77648 255134 77968 255218
rect 77648 254898 77690 255134
rect 77926 254898 77968 255134
rect 77648 254866 77968 254898
rect 108368 255454 108688 255486
rect 108368 255218 108410 255454
rect 108646 255218 108688 255454
rect 108368 255134 108688 255218
rect 108368 254898 108410 255134
rect 108646 254898 108688 255134
rect 108368 254866 108688 254898
rect 139088 255454 139408 255486
rect 139088 255218 139130 255454
rect 139366 255218 139408 255454
rect 139088 255134 139408 255218
rect 139088 254898 139130 255134
rect 139366 254898 139408 255134
rect 139088 254866 139408 254898
rect 169808 255454 170128 255486
rect 169808 255218 169850 255454
rect 170086 255218 170128 255454
rect 169808 255134 170128 255218
rect 169808 254898 169850 255134
rect 170086 254898 170128 255134
rect 169808 254866 170128 254898
rect 200528 255454 200848 255486
rect 200528 255218 200570 255454
rect 200806 255218 200848 255454
rect 200528 255134 200848 255218
rect 200528 254898 200570 255134
rect 200806 254898 200848 255134
rect 200528 254866 200848 254898
rect 231248 255454 231568 255486
rect 231248 255218 231290 255454
rect 231526 255218 231568 255454
rect 231248 255134 231568 255218
rect 231248 254898 231290 255134
rect 231526 254898 231568 255134
rect 231248 254866 231568 254898
rect 261968 255454 262288 255486
rect 261968 255218 262010 255454
rect 262246 255218 262288 255454
rect 261968 255134 262288 255218
rect 261968 254898 262010 255134
rect 262246 254898 262288 255134
rect 261968 254866 262288 254898
rect 292688 255454 293008 255486
rect 292688 255218 292730 255454
rect 292966 255218 293008 255454
rect 292688 255134 293008 255218
rect 292688 254898 292730 255134
rect 292966 254898 293008 255134
rect 292688 254866 293008 254898
rect 323408 255454 323728 255486
rect 323408 255218 323450 255454
rect 323686 255218 323728 255454
rect 323408 255134 323728 255218
rect 323408 254898 323450 255134
rect 323686 254898 323728 255134
rect 323408 254866 323728 254898
rect 354128 255454 354448 255486
rect 354128 255218 354170 255454
rect 354406 255218 354448 255454
rect 354128 255134 354448 255218
rect 354128 254898 354170 255134
rect 354406 254898 354448 255134
rect 354128 254866 354448 254898
rect 384848 255454 385168 255486
rect 384848 255218 384890 255454
rect 385126 255218 385168 255454
rect 384848 255134 385168 255218
rect 384848 254898 384890 255134
rect 385126 254898 385168 255134
rect 384848 254866 385168 254898
rect 415568 255454 415888 255486
rect 415568 255218 415610 255454
rect 415846 255218 415888 255454
rect 415568 255134 415888 255218
rect 415568 254898 415610 255134
rect 415846 254898 415888 255134
rect 415568 254866 415888 254898
rect 446288 255454 446608 255486
rect 446288 255218 446330 255454
rect 446566 255218 446608 255454
rect 446288 255134 446608 255218
rect 446288 254898 446330 255134
rect 446566 254898 446608 255134
rect 446288 254866 446608 254898
rect 477008 255454 477328 255486
rect 477008 255218 477050 255454
rect 477286 255218 477328 255454
rect 477008 255134 477328 255218
rect 477008 254898 477050 255134
rect 477286 254898 477328 255134
rect 477008 254866 477328 254898
rect 507728 255454 508048 255486
rect 507728 255218 507770 255454
rect 508006 255218 508048 255454
rect 507728 255134 508048 255218
rect 507728 254898 507770 255134
rect 508006 254898 508048 255134
rect 507728 254866 508048 254898
rect 538448 255454 538768 255486
rect 538448 255218 538490 255454
rect 538726 255218 538768 255454
rect 538448 255134 538768 255218
rect 538448 254898 538490 255134
rect 538726 254898 538768 255134
rect 538448 254866 538768 254898
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 31568 223174 31888 223206
rect 31568 222938 31610 223174
rect 31846 222938 31888 223174
rect 31568 222854 31888 222938
rect 31568 222618 31610 222854
rect 31846 222618 31888 222854
rect 31568 222586 31888 222618
rect 62288 223174 62608 223206
rect 62288 222938 62330 223174
rect 62566 222938 62608 223174
rect 62288 222854 62608 222938
rect 62288 222618 62330 222854
rect 62566 222618 62608 222854
rect 62288 222586 62608 222618
rect 93008 223174 93328 223206
rect 93008 222938 93050 223174
rect 93286 222938 93328 223174
rect 93008 222854 93328 222938
rect 93008 222618 93050 222854
rect 93286 222618 93328 222854
rect 93008 222586 93328 222618
rect 123728 223174 124048 223206
rect 123728 222938 123770 223174
rect 124006 222938 124048 223174
rect 123728 222854 124048 222938
rect 123728 222618 123770 222854
rect 124006 222618 124048 222854
rect 123728 222586 124048 222618
rect 154448 223174 154768 223206
rect 154448 222938 154490 223174
rect 154726 222938 154768 223174
rect 154448 222854 154768 222938
rect 154448 222618 154490 222854
rect 154726 222618 154768 222854
rect 154448 222586 154768 222618
rect 185168 223174 185488 223206
rect 185168 222938 185210 223174
rect 185446 222938 185488 223174
rect 185168 222854 185488 222938
rect 185168 222618 185210 222854
rect 185446 222618 185488 222854
rect 185168 222586 185488 222618
rect 215888 223174 216208 223206
rect 215888 222938 215930 223174
rect 216166 222938 216208 223174
rect 215888 222854 216208 222938
rect 215888 222618 215930 222854
rect 216166 222618 216208 222854
rect 215888 222586 216208 222618
rect 246608 223174 246928 223206
rect 246608 222938 246650 223174
rect 246886 222938 246928 223174
rect 246608 222854 246928 222938
rect 246608 222618 246650 222854
rect 246886 222618 246928 222854
rect 246608 222586 246928 222618
rect 277328 223174 277648 223206
rect 277328 222938 277370 223174
rect 277606 222938 277648 223174
rect 277328 222854 277648 222938
rect 277328 222618 277370 222854
rect 277606 222618 277648 222854
rect 277328 222586 277648 222618
rect 308048 223174 308368 223206
rect 308048 222938 308090 223174
rect 308326 222938 308368 223174
rect 308048 222854 308368 222938
rect 308048 222618 308090 222854
rect 308326 222618 308368 222854
rect 308048 222586 308368 222618
rect 338768 223174 339088 223206
rect 338768 222938 338810 223174
rect 339046 222938 339088 223174
rect 338768 222854 339088 222938
rect 338768 222618 338810 222854
rect 339046 222618 339088 222854
rect 338768 222586 339088 222618
rect 369488 223174 369808 223206
rect 369488 222938 369530 223174
rect 369766 222938 369808 223174
rect 369488 222854 369808 222938
rect 369488 222618 369530 222854
rect 369766 222618 369808 222854
rect 369488 222586 369808 222618
rect 400208 223174 400528 223206
rect 400208 222938 400250 223174
rect 400486 222938 400528 223174
rect 400208 222854 400528 222938
rect 400208 222618 400250 222854
rect 400486 222618 400528 222854
rect 400208 222586 400528 222618
rect 430928 223174 431248 223206
rect 430928 222938 430970 223174
rect 431206 222938 431248 223174
rect 430928 222854 431248 222938
rect 430928 222618 430970 222854
rect 431206 222618 431248 222854
rect 430928 222586 431248 222618
rect 461648 223174 461968 223206
rect 461648 222938 461690 223174
rect 461926 222938 461968 223174
rect 461648 222854 461968 222938
rect 461648 222618 461690 222854
rect 461926 222618 461968 222854
rect 461648 222586 461968 222618
rect 492368 223174 492688 223206
rect 492368 222938 492410 223174
rect 492646 222938 492688 223174
rect 492368 222854 492688 222938
rect 492368 222618 492410 222854
rect 492646 222618 492688 222854
rect 492368 222586 492688 222618
rect 523088 223174 523408 223206
rect 523088 222938 523130 223174
rect 523366 222938 523408 223174
rect 523088 222854 523408 222938
rect 523088 222618 523130 222854
rect 523366 222618 523408 222854
rect 523088 222586 523408 222618
rect 16208 219454 16528 219486
rect 16208 219218 16250 219454
rect 16486 219218 16528 219454
rect 16208 219134 16528 219218
rect 16208 218898 16250 219134
rect 16486 218898 16528 219134
rect 16208 218866 16528 218898
rect 46928 219454 47248 219486
rect 46928 219218 46970 219454
rect 47206 219218 47248 219454
rect 46928 219134 47248 219218
rect 46928 218898 46970 219134
rect 47206 218898 47248 219134
rect 46928 218866 47248 218898
rect 77648 219454 77968 219486
rect 77648 219218 77690 219454
rect 77926 219218 77968 219454
rect 77648 219134 77968 219218
rect 77648 218898 77690 219134
rect 77926 218898 77968 219134
rect 77648 218866 77968 218898
rect 108368 219454 108688 219486
rect 108368 219218 108410 219454
rect 108646 219218 108688 219454
rect 108368 219134 108688 219218
rect 108368 218898 108410 219134
rect 108646 218898 108688 219134
rect 108368 218866 108688 218898
rect 139088 219454 139408 219486
rect 139088 219218 139130 219454
rect 139366 219218 139408 219454
rect 139088 219134 139408 219218
rect 139088 218898 139130 219134
rect 139366 218898 139408 219134
rect 139088 218866 139408 218898
rect 169808 219454 170128 219486
rect 169808 219218 169850 219454
rect 170086 219218 170128 219454
rect 169808 219134 170128 219218
rect 169808 218898 169850 219134
rect 170086 218898 170128 219134
rect 169808 218866 170128 218898
rect 200528 219454 200848 219486
rect 200528 219218 200570 219454
rect 200806 219218 200848 219454
rect 200528 219134 200848 219218
rect 200528 218898 200570 219134
rect 200806 218898 200848 219134
rect 200528 218866 200848 218898
rect 231248 219454 231568 219486
rect 231248 219218 231290 219454
rect 231526 219218 231568 219454
rect 231248 219134 231568 219218
rect 231248 218898 231290 219134
rect 231526 218898 231568 219134
rect 231248 218866 231568 218898
rect 261968 219454 262288 219486
rect 261968 219218 262010 219454
rect 262246 219218 262288 219454
rect 261968 219134 262288 219218
rect 261968 218898 262010 219134
rect 262246 218898 262288 219134
rect 261968 218866 262288 218898
rect 292688 219454 293008 219486
rect 292688 219218 292730 219454
rect 292966 219218 293008 219454
rect 292688 219134 293008 219218
rect 292688 218898 292730 219134
rect 292966 218898 293008 219134
rect 292688 218866 293008 218898
rect 323408 219454 323728 219486
rect 323408 219218 323450 219454
rect 323686 219218 323728 219454
rect 323408 219134 323728 219218
rect 323408 218898 323450 219134
rect 323686 218898 323728 219134
rect 323408 218866 323728 218898
rect 354128 219454 354448 219486
rect 354128 219218 354170 219454
rect 354406 219218 354448 219454
rect 354128 219134 354448 219218
rect 354128 218898 354170 219134
rect 354406 218898 354448 219134
rect 354128 218866 354448 218898
rect 384848 219454 385168 219486
rect 384848 219218 384890 219454
rect 385126 219218 385168 219454
rect 384848 219134 385168 219218
rect 384848 218898 384890 219134
rect 385126 218898 385168 219134
rect 384848 218866 385168 218898
rect 415568 219454 415888 219486
rect 415568 219218 415610 219454
rect 415846 219218 415888 219454
rect 415568 219134 415888 219218
rect 415568 218898 415610 219134
rect 415846 218898 415888 219134
rect 415568 218866 415888 218898
rect 446288 219454 446608 219486
rect 446288 219218 446330 219454
rect 446566 219218 446608 219454
rect 446288 219134 446608 219218
rect 446288 218898 446330 219134
rect 446566 218898 446608 219134
rect 446288 218866 446608 218898
rect 477008 219454 477328 219486
rect 477008 219218 477050 219454
rect 477286 219218 477328 219454
rect 477008 219134 477328 219218
rect 477008 218898 477050 219134
rect 477286 218898 477328 219134
rect 477008 218866 477328 218898
rect 507728 219454 508048 219486
rect 507728 219218 507770 219454
rect 508006 219218 508048 219454
rect 507728 219134 508048 219218
rect 507728 218898 507770 219134
rect 508006 218898 508048 219134
rect 507728 218866 508048 218898
rect 538448 219454 538768 219486
rect 538448 219218 538490 219454
rect 538726 219218 538768 219454
rect 538448 219134 538768 219218
rect 538448 218898 538490 219134
rect 538726 218898 538768 219134
rect 538448 218866 538768 218898
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 31568 187174 31888 187206
rect 31568 186938 31610 187174
rect 31846 186938 31888 187174
rect 31568 186854 31888 186938
rect 31568 186618 31610 186854
rect 31846 186618 31888 186854
rect 31568 186586 31888 186618
rect 62288 187174 62608 187206
rect 62288 186938 62330 187174
rect 62566 186938 62608 187174
rect 62288 186854 62608 186938
rect 62288 186618 62330 186854
rect 62566 186618 62608 186854
rect 62288 186586 62608 186618
rect 93008 187174 93328 187206
rect 93008 186938 93050 187174
rect 93286 186938 93328 187174
rect 93008 186854 93328 186938
rect 93008 186618 93050 186854
rect 93286 186618 93328 186854
rect 93008 186586 93328 186618
rect 123728 187174 124048 187206
rect 123728 186938 123770 187174
rect 124006 186938 124048 187174
rect 123728 186854 124048 186938
rect 123728 186618 123770 186854
rect 124006 186618 124048 186854
rect 123728 186586 124048 186618
rect 154448 187174 154768 187206
rect 154448 186938 154490 187174
rect 154726 186938 154768 187174
rect 154448 186854 154768 186938
rect 154448 186618 154490 186854
rect 154726 186618 154768 186854
rect 154448 186586 154768 186618
rect 185168 187174 185488 187206
rect 185168 186938 185210 187174
rect 185446 186938 185488 187174
rect 185168 186854 185488 186938
rect 185168 186618 185210 186854
rect 185446 186618 185488 186854
rect 185168 186586 185488 186618
rect 215888 187174 216208 187206
rect 215888 186938 215930 187174
rect 216166 186938 216208 187174
rect 215888 186854 216208 186938
rect 215888 186618 215930 186854
rect 216166 186618 216208 186854
rect 215888 186586 216208 186618
rect 246608 187174 246928 187206
rect 246608 186938 246650 187174
rect 246886 186938 246928 187174
rect 246608 186854 246928 186938
rect 246608 186618 246650 186854
rect 246886 186618 246928 186854
rect 246608 186586 246928 186618
rect 277328 187174 277648 187206
rect 277328 186938 277370 187174
rect 277606 186938 277648 187174
rect 277328 186854 277648 186938
rect 277328 186618 277370 186854
rect 277606 186618 277648 186854
rect 277328 186586 277648 186618
rect 308048 187174 308368 187206
rect 308048 186938 308090 187174
rect 308326 186938 308368 187174
rect 308048 186854 308368 186938
rect 308048 186618 308090 186854
rect 308326 186618 308368 186854
rect 308048 186586 308368 186618
rect 338768 187174 339088 187206
rect 338768 186938 338810 187174
rect 339046 186938 339088 187174
rect 338768 186854 339088 186938
rect 338768 186618 338810 186854
rect 339046 186618 339088 186854
rect 338768 186586 339088 186618
rect 369488 187174 369808 187206
rect 369488 186938 369530 187174
rect 369766 186938 369808 187174
rect 369488 186854 369808 186938
rect 369488 186618 369530 186854
rect 369766 186618 369808 186854
rect 369488 186586 369808 186618
rect 400208 187174 400528 187206
rect 400208 186938 400250 187174
rect 400486 186938 400528 187174
rect 400208 186854 400528 186938
rect 400208 186618 400250 186854
rect 400486 186618 400528 186854
rect 400208 186586 400528 186618
rect 430928 187174 431248 187206
rect 430928 186938 430970 187174
rect 431206 186938 431248 187174
rect 430928 186854 431248 186938
rect 430928 186618 430970 186854
rect 431206 186618 431248 186854
rect 430928 186586 431248 186618
rect 461648 187174 461968 187206
rect 461648 186938 461690 187174
rect 461926 186938 461968 187174
rect 461648 186854 461968 186938
rect 461648 186618 461690 186854
rect 461926 186618 461968 186854
rect 461648 186586 461968 186618
rect 492368 187174 492688 187206
rect 492368 186938 492410 187174
rect 492646 186938 492688 187174
rect 492368 186854 492688 186938
rect 492368 186618 492410 186854
rect 492646 186618 492688 186854
rect 492368 186586 492688 186618
rect 523088 187174 523408 187206
rect 523088 186938 523130 187174
rect 523366 186938 523408 187174
rect 523088 186854 523408 186938
rect 523088 186618 523130 186854
rect 523366 186618 523408 186854
rect 523088 186586 523408 186618
rect 16208 183454 16528 183486
rect 16208 183218 16250 183454
rect 16486 183218 16528 183454
rect 16208 183134 16528 183218
rect 16208 182898 16250 183134
rect 16486 182898 16528 183134
rect 16208 182866 16528 182898
rect 46928 183454 47248 183486
rect 46928 183218 46970 183454
rect 47206 183218 47248 183454
rect 46928 183134 47248 183218
rect 46928 182898 46970 183134
rect 47206 182898 47248 183134
rect 46928 182866 47248 182898
rect 77648 183454 77968 183486
rect 77648 183218 77690 183454
rect 77926 183218 77968 183454
rect 77648 183134 77968 183218
rect 77648 182898 77690 183134
rect 77926 182898 77968 183134
rect 77648 182866 77968 182898
rect 108368 183454 108688 183486
rect 108368 183218 108410 183454
rect 108646 183218 108688 183454
rect 108368 183134 108688 183218
rect 108368 182898 108410 183134
rect 108646 182898 108688 183134
rect 108368 182866 108688 182898
rect 139088 183454 139408 183486
rect 139088 183218 139130 183454
rect 139366 183218 139408 183454
rect 139088 183134 139408 183218
rect 139088 182898 139130 183134
rect 139366 182898 139408 183134
rect 139088 182866 139408 182898
rect 169808 183454 170128 183486
rect 169808 183218 169850 183454
rect 170086 183218 170128 183454
rect 169808 183134 170128 183218
rect 169808 182898 169850 183134
rect 170086 182898 170128 183134
rect 169808 182866 170128 182898
rect 200528 183454 200848 183486
rect 200528 183218 200570 183454
rect 200806 183218 200848 183454
rect 200528 183134 200848 183218
rect 200528 182898 200570 183134
rect 200806 182898 200848 183134
rect 200528 182866 200848 182898
rect 231248 183454 231568 183486
rect 231248 183218 231290 183454
rect 231526 183218 231568 183454
rect 231248 183134 231568 183218
rect 231248 182898 231290 183134
rect 231526 182898 231568 183134
rect 231248 182866 231568 182898
rect 261968 183454 262288 183486
rect 261968 183218 262010 183454
rect 262246 183218 262288 183454
rect 261968 183134 262288 183218
rect 261968 182898 262010 183134
rect 262246 182898 262288 183134
rect 261968 182866 262288 182898
rect 292688 183454 293008 183486
rect 292688 183218 292730 183454
rect 292966 183218 293008 183454
rect 292688 183134 293008 183218
rect 292688 182898 292730 183134
rect 292966 182898 293008 183134
rect 292688 182866 293008 182898
rect 323408 183454 323728 183486
rect 323408 183218 323450 183454
rect 323686 183218 323728 183454
rect 323408 183134 323728 183218
rect 323408 182898 323450 183134
rect 323686 182898 323728 183134
rect 323408 182866 323728 182898
rect 354128 183454 354448 183486
rect 354128 183218 354170 183454
rect 354406 183218 354448 183454
rect 354128 183134 354448 183218
rect 354128 182898 354170 183134
rect 354406 182898 354448 183134
rect 354128 182866 354448 182898
rect 384848 183454 385168 183486
rect 384848 183218 384890 183454
rect 385126 183218 385168 183454
rect 384848 183134 385168 183218
rect 384848 182898 384890 183134
rect 385126 182898 385168 183134
rect 384848 182866 385168 182898
rect 415568 183454 415888 183486
rect 415568 183218 415610 183454
rect 415846 183218 415888 183454
rect 415568 183134 415888 183218
rect 415568 182898 415610 183134
rect 415846 182898 415888 183134
rect 415568 182866 415888 182898
rect 446288 183454 446608 183486
rect 446288 183218 446330 183454
rect 446566 183218 446608 183454
rect 446288 183134 446608 183218
rect 446288 182898 446330 183134
rect 446566 182898 446608 183134
rect 446288 182866 446608 182898
rect 477008 183454 477328 183486
rect 477008 183218 477050 183454
rect 477286 183218 477328 183454
rect 477008 183134 477328 183218
rect 477008 182898 477050 183134
rect 477286 182898 477328 183134
rect 477008 182866 477328 182898
rect 507728 183454 508048 183486
rect 507728 183218 507770 183454
rect 508006 183218 508048 183454
rect 507728 183134 508048 183218
rect 507728 182898 507770 183134
rect 508006 182898 508048 183134
rect 507728 182866 508048 182898
rect 538448 183454 538768 183486
rect 538448 183218 538490 183454
rect 538726 183218 538768 183454
rect 538448 183134 538768 183218
rect 538448 182898 538490 183134
rect 538726 182898 538768 183134
rect 538448 182866 538768 182898
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 31568 151174 31888 151206
rect 31568 150938 31610 151174
rect 31846 150938 31888 151174
rect 31568 150854 31888 150938
rect 31568 150618 31610 150854
rect 31846 150618 31888 150854
rect 31568 150586 31888 150618
rect 62288 151174 62608 151206
rect 62288 150938 62330 151174
rect 62566 150938 62608 151174
rect 62288 150854 62608 150938
rect 62288 150618 62330 150854
rect 62566 150618 62608 150854
rect 62288 150586 62608 150618
rect 93008 151174 93328 151206
rect 93008 150938 93050 151174
rect 93286 150938 93328 151174
rect 93008 150854 93328 150938
rect 93008 150618 93050 150854
rect 93286 150618 93328 150854
rect 93008 150586 93328 150618
rect 123728 151174 124048 151206
rect 123728 150938 123770 151174
rect 124006 150938 124048 151174
rect 123728 150854 124048 150938
rect 123728 150618 123770 150854
rect 124006 150618 124048 150854
rect 123728 150586 124048 150618
rect 154448 151174 154768 151206
rect 154448 150938 154490 151174
rect 154726 150938 154768 151174
rect 154448 150854 154768 150938
rect 154448 150618 154490 150854
rect 154726 150618 154768 150854
rect 154448 150586 154768 150618
rect 185168 151174 185488 151206
rect 185168 150938 185210 151174
rect 185446 150938 185488 151174
rect 185168 150854 185488 150938
rect 185168 150618 185210 150854
rect 185446 150618 185488 150854
rect 185168 150586 185488 150618
rect 215888 151174 216208 151206
rect 215888 150938 215930 151174
rect 216166 150938 216208 151174
rect 215888 150854 216208 150938
rect 215888 150618 215930 150854
rect 216166 150618 216208 150854
rect 215888 150586 216208 150618
rect 246608 151174 246928 151206
rect 246608 150938 246650 151174
rect 246886 150938 246928 151174
rect 246608 150854 246928 150938
rect 246608 150618 246650 150854
rect 246886 150618 246928 150854
rect 246608 150586 246928 150618
rect 277328 151174 277648 151206
rect 277328 150938 277370 151174
rect 277606 150938 277648 151174
rect 277328 150854 277648 150938
rect 277328 150618 277370 150854
rect 277606 150618 277648 150854
rect 277328 150586 277648 150618
rect 308048 151174 308368 151206
rect 308048 150938 308090 151174
rect 308326 150938 308368 151174
rect 308048 150854 308368 150938
rect 308048 150618 308090 150854
rect 308326 150618 308368 150854
rect 308048 150586 308368 150618
rect 338768 151174 339088 151206
rect 338768 150938 338810 151174
rect 339046 150938 339088 151174
rect 338768 150854 339088 150938
rect 338768 150618 338810 150854
rect 339046 150618 339088 150854
rect 338768 150586 339088 150618
rect 369488 151174 369808 151206
rect 369488 150938 369530 151174
rect 369766 150938 369808 151174
rect 369488 150854 369808 150938
rect 369488 150618 369530 150854
rect 369766 150618 369808 150854
rect 369488 150586 369808 150618
rect 400208 151174 400528 151206
rect 400208 150938 400250 151174
rect 400486 150938 400528 151174
rect 400208 150854 400528 150938
rect 400208 150618 400250 150854
rect 400486 150618 400528 150854
rect 400208 150586 400528 150618
rect 430928 151174 431248 151206
rect 430928 150938 430970 151174
rect 431206 150938 431248 151174
rect 430928 150854 431248 150938
rect 430928 150618 430970 150854
rect 431206 150618 431248 150854
rect 430928 150586 431248 150618
rect 461648 151174 461968 151206
rect 461648 150938 461690 151174
rect 461926 150938 461968 151174
rect 461648 150854 461968 150938
rect 461648 150618 461690 150854
rect 461926 150618 461968 150854
rect 461648 150586 461968 150618
rect 492368 151174 492688 151206
rect 492368 150938 492410 151174
rect 492646 150938 492688 151174
rect 492368 150854 492688 150938
rect 492368 150618 492410 150854
rect 492646 150618 492688 150854
rect 492368 150586 492688 150618
rect 523088 151174 523408 151206
rect 523088 150938 523130 151174
rect 523366 150938 523408 151174
rect 523088 150854 523408 150938
rect 523088 150618 523130 150854
rect 523366 150618 523408 150854
rect 523088 150586 523408 150618
rect 16208 147454 16528 147486
rect 16208 147218 16250 147454
rect 16486 147218 16528 147454
rect 16208 147134 16528 147218
rect 16208 146898 16250 147134
rect 16486 146898 16528 147134
rect 16208 146866 16528 146898
rect 46928 147454 47248 147486
rect 46928 147218 46970 147454
rect 47206 147218 47248 147454
rect 46928 147134 47248 147218
rect 46928 146898 46970 147134
rect 47206 146898 47248 147134
rect 46928 146866 47248 146898
rect 77648 147454 77968 147486
rect 77648 147218 77690 147454
rect 77926 147218 77968 147454
rect 77648 147134 77968 147218
rect 77648 146898 77690 147134
rect 77926 146898 77968 147134
rect 77648 146866 77968 146898
rect 108368 147454 108688 147486
rect 108368 147218 108410 147454
rect 108646 147218 108688 147454
rect 108368 147134 108688 147218
rect 108368 146898 108410 147134
rect 108646 146898 108688 147134
rect 108368 146866 108688 146898
rect 139088 147454 139408 147486
rect 139088 147218 139130 147454
rect 139366 147218 139408 147454
rect 139088 147134 139408 147218
rect 139088 146898 139130 147134
rect 139366 146898 139408 147134
rect 139088 146866 139408 146898
rect 169808 147454 170128 147486
rect 169808 147218 169850 147454
rect 170086 147218 170128 147454
rect 169808 147134 170128 147218
rect 169808 146898 169850 147134
rect 170086 146898 170128 147134
rect 169808 146866 170128 146898
rect 200528 147454 200848 147486
rect 200528 147218 200570 147454
rect 200806 147218 200848 147454
rect 200528 147134 200848 147218
rect 200528 146898 200570 147134
rect 200806 146898 200848 147134
rect 200528 146866 200848 146898
rect 231248 147454 231568 147486
rect 231248 147218 231290 147454
rect 231526 147218 231568 147454
rect 231248 147134 231568 147218
rect 231248 146898 231290 147134
rect 231526 146898 231568 147134
rect 231248 146866 231568 146898
rect 261968 147454 262288 147486
rect 261968 147218 262010 147454
rect 262246 147218 262288 147454
rect 261968 147134 262288 147218
rect 261968 146898 262010 147134
rect 262246 146898 262288 147134
rect 261968 146866 262288 146898
rect 292688 147454 293008 147486
rect 292688 147218 292730 147454
rect 292966 147218 293008 147454
rect 292688 147134 293008 147218
rect 292688 146898 292730 147134
rect 292966 146898 293008 147134
rect 292688 146866 293008 146898
rect 323408 147454 323728 147486
rect 323408 147218 323450 147454
rect 323686 147218 323728 147454
rect 323408 147134 323728 147218
rect 323408 146898 323450 147134
rect 323686 146898 323728 147134
rect 323408 146866 323728 146898
rect 354128 147454 354448 147486
rect 354128 147218 354170 147454
rect 354406 147218 354448 147454
rect 354128 147134 354448 147218
rect 354128 146898 354170 147134
rect 354406 146898 354448 147134
rect 354128 146866 354448 146898
rect 384848 147454 385168 147486
rect 384848 147218 384890 147454
rect 385126 147218 385168 147454
rect 384848 147134 385168 147218
rect 384848 146898 384890 147134
rect 385126 146898 385168 147134
rect 384848 146866 385168 146898
rect 415568 147454 415888 147486
rect 415568 147218 415610 147454
rect 415846 147218 415888 147454
rect 415568 147134 415888 147218
rect 415568 146898 415610 147134
rect 415846 146898 415888 147134
rect 415568 146866 415888 146898
rect 446288 147454 446608 147486
rect 446288 147218 446330 147454
rect 446566 147218 446608 147454
rect 446288 147134 446608 147218
rect 446288 146898 446330 147134
rect 446566 146898 446608 147134
rect 446288 146866 446608 146898
rect 477008 147454 477328 147486
rect 477008 147218 477050 147454
rect 477286 147218 477328 147454
rect 477008 147134 477328 147218
rect 477008 146898 477050 147134
rect 477286 146898 477328 147134
rect 477008 146866 477328 146898
rect 507728 147454 508048 147486
rect 507728 147218 507770 147454
rect 508006 147218 508048 147454
rect 507728 147134 508048 147218
rect 507728 146898 507770 147134
rect 508006 146898 508048 147134
rect 507728 146866 508048 146898
rect 538448 147454 538768 147486
rect 538448 147218 538490 147454
rect 538726 147218 538768 147454
rect 538448 147134 538768 147218
rect 538448 146898 538490 147134
rect 538726 146898 538768 147134
rect 538448 146866 538768 146898
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 31568 115174 31888 115206
rect 31568 114938 31610 115174
rect 31846 114938 31888 115174
rect 31568 114854 31888 114938
rect 31568 114618 31610 114854
rect 31846 114618 31888 114854
rect 31568 114586 31888 114618
rect 62288 115174 62608 115206
rect 62288 114938 62330 115174
rect 62566 114938 62608 115174
rect 62288 114854 62608 114938
rect 62288 114618 62330 114854
rect 62566 114618 62608 114854
rect 62288 114586 62608 114618
rect 93008 115174 93328 115206
rect 93008 114938 93050 115174
rect 93286 114938 93328 115174
rect 93008 114854 93328 114938
rect 93008 114618 93050 114854
rect 93286 114618 93328 114854
rect 93008 114586 93328 114618
rect 123728 115174 124048 115206
rect 123728 114938 123770 115174
rect 124006 114938 124048 115174
rect 123728 114854 124048 114938
rect 123728 114618 123770 114854
rect 124006 114618 124048 114854
rect 123728 114586 124048 114618
rect 154448 115174 154768 115206
rect 154448 114938 154490 115174
rect 154726 114938 154768 115174
rect 154448 114854 154768 114938
rect 154448 114618 154490 114854
rect 154726 114618 154768 114854
rect 154448 114586 154768 114618
rect 185168 115174 185488 115206
rect 185168 114938 185210 115174
rect 185446 114938 185488 115174
rect 185168 114854 185488 114938
rect 185168 114618 185210 114854
rect 185446 114618 185488 114854
rect 185168 114586 185488 114618
rect 215888 115174 216208 115206
rect 215888 114938 215930 115174
rect 216166 114938 216208 115174
rect 215888 114854 216208 114938
rect 215888 114618 215930 114854
rect 216166 114618 216208 114854
rect 215888 114586 216208 114618
rect 246608 115174 246928 115206
rect 246608 114938 246650 115174
rect 246886 114938 246928 115174
rect 246608 114854 246928 114938
rect 246608 114618 246650 114854
rect 246886 114618 246928 114854
rect 246608 114586 246928 114618
rect 277328 115174 277648 115206
rect 277328 114938 277370 115174
rect 277606 114938 277648 115174
rect 277328 114854 277648 114938
rect 277328 114618 277370 114854
rect 277606 114618 277648 114854
rect 277328 114586 277648 114618
rect 308048 115174 308368 115206
rect 308048 114938 308090 115174
rect 308326 114938 308368 115174
rect 308048 114854 308368 114938
rect 308048 114618 308090 114854
rect 308326 114618 308368 114854
rect 308048 114586 308368 114618
rect 338768 115174 339088 115206
rect 338768 114938 338810 115174
rect 339046 114938 339088 115174
rect 338768 114854 339088 114938
rect 338768 114618 338810 114854
rect 339046 114618 339088 114854
rect 338768 114586 339088 114618
rect 369488 115174 369808 115206
rect 369488 114938 369530 115174
rect 369766 114938 369808 115174
rect 369488 114854 369808 114938
rect 369488 114618 369530 114854
rect 369766 114618 369808 114854
rect 369488 114586 369808 114618
rect 400208 115174 400528 115206
rect 400208 114938 400250 115174
rect 400486 114938 400528 115174
rect 400208 114854 400528 114938
rect 400208 114618 400250 114854
rect 400486 114618 400528 114854
rect 400208 114586 400528 114618
rect 430928 115174 431248 115206
rect 430928 114938 430970 115174
rect 431206 114938 431248 115174
rect 430928 114854 431248 114938
rect 430928 114618 430970 114854
rect 431206 114618 431248 114854
rect 430928 114586 431248 114618
rect 461648 115174 461968 115206
rect 461648 114938 461690 115174
rect 461926 114938 461968 115174
rect 461648 114854 461968 114938
rect 461648 114618 461690 114854
rect 461926 114618 461968 114854
rect 461648 114586 461968 114618
rect 492368 115174 492688 115206
rect 492368 114938 492410 115174
rect 492646 114938 492688 115174
rect 492368 114854 492688 114938
rect 492368 114618 492410 114854
rect 492646 114618 492688 114854
rect 492368 114586 492688 114618
rect 523088 115174 523408 115206
rect 523088 114938 523130 115174
rect 523366 114938 523408 115174
rect 523088 114854 523408 114938
rect 523088 114618 523130 114854
rect 523366 114618 523408 114854
rect 523088 114586 523408 114618
rect 16208 111454 16528 111486
rect 16208 111218 16250 111454
rect 16486 111218 16528 111454
rect 16208 111134 16528 111218
rect 16208 110898 16250 111134
rect 16486 110898 16528 111134
rect 16208 110866 16528 110898
rect 46928 111454 47248 111486
rect 46928 111218 46970 111454
rect 47206 111218 47248 111454
rect 46928 111134 47248 111218
rect 46928 110898 46970 111134
rect 47206 110898 47248 111134
rect 46928 110866 47248 110898
rect 77648 111454 77968 111486
rect 77648 111218 77690 111454
rect 77926 111218 77968 111454
rect 77648 111134 77968 111218
rect 77648 110898 77690 111134
rect 77926 110898 77968 111134
rect 77648 110866 77968 110898
rect 108368 111454 108688 111486
rect 108368 111218 108410 111454
rect 108646 111218 108688 111454
rect 108368 111134 108688 111218
rect 108368 110898 108410 111134
rect 108646 110898 108688 111134
rect 108368 110866 108688 110898
rect 139088 111454 139408 111486
rect 139088 111218 139130 111454
rect 139366 111218 139408 111454
rect 139088 111134 139408 111218
rect 139088 110898 139130 111134
rect 139366 110898 139408 111134
rect 139088 110866 139408 110898
rect 169808 111454 170128 111486
rect 169808 111218 169850 111454
rect 170086 111218 170128 111454
rect 169808 111134 170128 111218
rect 169808 110898 169850 111134
rect 170086 110898 170128 111134
rect 169808 110866 170128 110898
rect 200528 111454 200848 111486
rect 200528 111218 200570 111454
rect 200806 111218 200848 111454
rect 200528 111134 200848 111218
rect 200528 110898 200570 111134
rect 200806 110898 200848 111134
rect 200528 110866 200848 110898
rect 231248 111454 231568 111486
rect 231248 111218 231290 111454
rect 231526 111218 231568 111454
rect 231248 111134 231568 111218
rect 231248 110898 231290 111134
rect 231526 110898 231568 111134
rect 231248 110866 231568 110898
rect 261968 111454 262288 111486
rect 261968 111218 262010 111454
rect 262246 111218 262288 111454
rect 261968 111134 262288 111218
rect 261968 110898 262010 111134
rect 262246 110898 262288 111134
rect 261968 110866 262288 110898
rect 292688 111454 293008 111486
rect 292688 111218 292730 111454
rect 292966 111218 293008 111454
rect 292688 111134 293008 111218
rect 292688 110898 292730 111134
rect 292966 110898 293008 111134
rect 292688 110866 293008 110898
rect 323408 111454 323728 111486
rect 323408 111218 323450 111454
rect 323686 111218 323728 111454
rect 323408 111134 323728 111218
rect 323408 110898 323450 111134
rect 323686 110898 323728 111134
rect 323408 110866 323728 110898
rect 354128 111454 354448 111486
rect 354128 111218 354170 111454
rect 354406 111218 354448 111454
rect 354128 111134 354448 111218
rect 354128 110898 354170 111134
rect 354406 110898 354448 111134
rect 354128 110866 354448 110898
rect 384848 111454 385168 111486
rect 384848 111218 384890 111454
rect 385126 111218 385168 111454
rect 384848 111134 385168 111218
rect 384848 110898 384890 111134
rect 385126 110898 385168 111134
rect 384848 110866 385168 110898
rect 415568 111454 415888 111486
rect 415568 111218 415610 111454
rect 415846 111218 415888 111454
rect 415568 111134 415888 111218
rect 415568 110898 415610 111134
rect 415846 110898 415888 111134
rect 415568 110866 415888 110898
rect 446288 111454 446608 111486
rect 446288 111218 446330 111454
rect 446566 111218 446608 111454
rect 446288 111134 446608 111218
rect 446288 110898 446330 111134
rect 446566 110898 446608 111134
rect 446288 110866 446608 110898
rect 477008 111454 477328 111486
rect 477008 111218 477050 111454
rect 477286 111218 477328 111454
rect 477008 111134 477328 111218
rect 477008 110898 477050 111134
rect 477286 110898 477328 111134
rect 477008 110866 477328 110898
rect 507728 111454 508048 111486
rect 507728 111218 507770 111454
rect 508006 111218 508048 111454
rect 507728 111134 508048 111218
rect 507728 110898 507770 111134
rect 508006 110898 508048 111134
rect 507728 110866 508048 110898
rect 538448 111454 538768 111486
rect 538448 111218 538490 111454
rect 538726 111218 538768 111454
rect 538448 111134 538768 111218
rect 538448 110898 538490 111134
rect 538726 110898 538768 111134
rect 538448 110866 538768 110898
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 31568 79174 31888 79206
rect 31568 78938 31610 79174
rect 31846 78938 31888 79174
rect 31568 78854 31888 78938
rect 31568 78618 31610 78854
rect 31846 78618 31888 78854
rect 31568 78586 31888 78618
rect 62288 79174 62608 79206
rect 62288 78938 62330 79174
rect 62566 78938 62608 79174
rect 62288 78854 62608 78938
rect 62288 78618 62330 78854
rect 62566 78618 62608 78854
rect 62288 78586 62608 78618
rect 93008 79174 93328 79206
rect 93008 78938 93050 79174
rect 93286 78938 93328 79174
rect 93008 78854 93328 78938
rect 93008 78618 93050 78854
rect 93286 78618 93328 78854
rect 93008 78586 93328 78618
rect 123728 79174 124048 79206
rect 123728 78938 123770 79174
rect 124006 78938 124048 79174
rect 123728 78854 124048 78938
rect 123728 78618 123770 78854
rect 124006 78618 124048 78854
rect 123728 78586 124048 78618
rect 154448 79174 154768 79206
rect 154448 78938 154490 79174
rect 154726 78938 154768 79174
rect 154448 78854 154768 78938
rect 154448 78618 154490 78854
rect 154726 78618 154768 78854
rect 154448 78586 154768 78618
rect 185168 79174 185488 79206
rect 185168 78938 185210 79174
rect 185446 78938 185488 79174
rect 185168 78854 185488 78938
rect 185168 78618 185210 78854
rect 185446 78618 185488 78854
rect 185168 78586 185488 78618
rect 215888 79174 216208 79206
rect 215888 78938 215930 79174
rect 216166 78938 216208 79174
rect 215888 78854 216208 78938
rect 215888 78618 215930 78854
rect 216166 78618 216208 78854
rect 215888 78586 216208 78618
rect 246608 79174 246928 79206
rect 246608 78938 246650 79174
rect 246886 78938 246928 79174
rect 246608 78854 246928 78938
rect 246608 78618 246650 78854
rect 246886 78618 246928 78854
rect 246608 78586 246928 78618
rect 277328 79174 277648 79206
rect 277328 78938 277370 79174
rect 277606 78938 277648 79174
rect 277328 78854 277648 78938
rect 277328 78618 277370 78854
rect 277606 78618 277648 78854
rect 277328 78586 277648 78618
rect 308048 79174 308368 79206
rect 308048 78938 308090 79174
rect 308326 78938 308368 79174
rect 308048 78854 308368 78938
rect 308048 78618 308090 78854
rect 308326 78618 308368 78854
rect 308048 78586 308368 78618
rect 338768 79174 339088 79206
rect 338768 78938 338810 79174
rect 339046 78938 339088 79174
rect 338768 78854 339088 78938
rect 338768 78618 338810 78854
rect 339046 78618 339088 78854
rect 338768 78586 339088 78618
rect 369488 79174 369808 79206
rect 369488 78938 369530 79174
rect 369766 78938 369808 79174
rect 369488 78854 369808 78938
rect 369488 78618 369530 78854
rect 369766 78618 369808 78854
rect 369488 78586 369808 78618
rect 400208 79174 400528 79206
rect 400208 78938 400250 79174
rect 400486 78938 400528 79174
rect 400208 78854 400528 78938
rect 400208 78618 400250 78854
rect 400486 78618 400528 78854
rect 400208 78586 400528 78618
rect 430928 79174 431248 79206
rect 430928 78938 430970 79174
rect 431206 78938 431248 79174
rect 430928 78854 431248 78938
rect 430928 78618 430970 78854
rect 431206 78618 431248 78854
rect 430928 78586 431248 78618
rect 461648 79174 461968 79206
rect 461648 78938 461690 79174
rect 461926 78938 461968 79174
rect 461648 78854 461968 78938
rect 461648 78618 461690 78854
rect 461926 78618 461968 78854
rect 461648 78586 461968 78618
rect 492368 79174 492688 79206
rect 492368 78938 492410 79174
rect 492646 78938 492688 79174
rect 492368 78854 492688 78938
rect 492368 78618 492410 78854
rect 492646 78618 492688 78854
rect 492368 78586 492688 78618
rect 523088 79174 523408 79206
rect 523088 78938 523130 79174
rect 523366 78938 523408 79174
rect 523088 78854 523408 78938
rect 523088 78618 523130 78854
rect 523366 78618 523408 78854
rect 523088 78586 523408 78618
rect 16208 75454 16528 75486
rect 16208 75218 16250 75454
rect 16486 75218 16528 75454
rect 16208 75134 16528 75218
rect 16208 74898 16250 75134
rect 16486 74898 16528 75134
rect 16208 74866 16528 74898
rect 46928 75454 47248 75486
rect 46928 75218 46970 75454
rect 47206 75218 47248 75454
rect 46928 75134 47248 75218
rect 46928 74898 46970 75134
rect 47206 74898 47248 75134
rect 46928 74866 47248 74898
rect 77648 75454 77968 75486
rect 77648 75218 77690 75454
rect 77926 75218 77968 75454
rect 77648 75134 77968 75218
rect 77648 74898 77690 75134
rect 77926 74898 77968 75134
rect 77648 74866 77968 74898
rect 108368 75454 108688 75486
rect 108368 75218 108410 75454
rect 108646 75218 108688 75454
rect 108368 75134 108688 75218
rect 108368 74898 108410 75134
rect 108646 74898 108688 75134
rect 108368 74866 108688 74898
rect 139088 75454 139408 75486
rect 139088 75218 139130 75454
rect 139366 75218 139408 75454
rect 139088 75134 139408 75218
rect 139088 74898 139130 75134
rect 139366 74898 139408 75134
rect 139088 74866 139408 74898
rect 169808 75454 170128 75486
rect 169808 75218 169850 75454
rect 170086 75218 170128 75454
rect 169808 75134 170128 75218
rect 169808 74898 169850 75134
rect 170086 74898 170128 75134
rect 169808 74866 170128 74898
rect 200528 75454 200848 75486
rect 200528 75218 200570 75454
rect 200806 75218 200848 75454
rect 200528 75134 200848 75218
rect 200528 74898 200570 75134
rect 200806 74898 200848 75134
rect 200528 74866 200848 74898
rect 231248 75454 231568 75486
rect 231248 75218 231290 75454
rect 231526 75218 231568 75454
rect 231248 75134 231568 75218
rect 231248 74898 231290 75134
rect 231526 74898 231568 75134
rect 231248 74866 231568 74898
rect 261968 75454 262288 75486
rect 261968 75218 262010 75454
rect 262246 75218 262288 75454
rect 261968 75134 262288 75218
rect 261968 74898 262010 75134
rect 262246 74898 262288 75134
rect 261968 74866 262288 74898
rect 292688 75454 293008 75486
rect 292688 75218 292730 75454
rect 292966 75218 293008 75454
rect 292688 75134 293008 75218
rect 292688 74898 292730 75134
rect 292966 74898 293008 75134
rect 292688 74866 293008 74898
rect 323408 75454 323728 75486
rect 323408 75218 323450 75454
rect 323686 75218 323728 75454
rect 323408 75134 323728 75218
rect 323408 74898 323450 75134
rect 323686 74898 323728 75134
rect 323408 74866 323728 74898
rect 354128 75454 354448 75486
rect 354128 75218 354170 75454
rect 354406 75218 354448 75454
rect 354128 75134 354448 75218
rect 354128 74898 354170 75134
rect 354406 74898 354448 75134
rect 354128 74866 354448 74898
rect 384848 75454 385168 75486
rect 384848 75218 384890 75454
rect 385126 75218 385168 75454
rect 384848 75134 385168 75218
rect 384848 74898 384890 75134
rect 385126 74898 385168 75134
rect 384848 74866 385168 74898
rect 415568 75454 415888 75486
rect 415568 75218 415610 75454
rect 415846 75218 415888 75454
rect 415568 75134 415888 75218
rect 415568 74898 415610 75134
rect 415846 74898 415888 75134
rect 415568 74866 415888 74898
rect 446288 75454 446608 75486
rect 446288 75218 446330 75454
rect 446566 75218 446608 75454
rect 446288 75134 446608 75218
rect 446288 74898 446330 75134
rect 446566 74898 446608 75134
rect 446288 74866 446608 74898
rect 477008 75454 477328 75486
rect 477008 75218 477050 75454
rect 477286 75218 477328 75454
rect 477008 75134 477328 75218
rect 477008 74898 477050 75134
rect 477286 74898 477328 75134
rect 477008 74866 477328 74898
rect 507728 75454 508048 75486
rect 507728 75218 507770 75454
rect 508006 75218 508048 75454
rect 507728 75134 508048 75218
rect 507728 74898 507770 75134
rect 508006 74898 508048 75134
rect 507728 74866 508048 74898
rect 538448 75454 538768 75486
rect 538448 75218 538490 75454
rect 538726 75218 538768 75454
rect 538448 75134 538768 75218
rect 538448 74898 538490 75134
rect 538726 74898 538768 75134
rect 538448 74866 538768 74898
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 31568 43174 31888 43206
rect 31568 42938 31610 43174
rect 31846 42938 31888 43174
rect 31568 42854 31888 42938
rect 31568 42618 31610 42854
rect 31846 42618 31888 42854
rect 31568 42586 31888 42618
rect 62288 43174 62608 43206
rect 62288 42938 62330 43174
rect 62566 42938 62608 43174
rect 62288 42854 62608 42938
rect 62288 42618 62330 42854
rect 62566 42618 62608 42854
rect 62288 42586 62608 42618
rect 93008 43174 93328 43206
rect 93008 42938 93050 43174
rect 93286 42938 93328 43174
rect 93008 42854 93328 42938
rect 93008 42618 93050 42854
rect 93286 42618 93328 42854
rect 93008 42586 93328 42618
rect 123728 43174 124048 43206
rect 123728 42938 123770 43174
rect 124006 42938 124048 43174
rect 123728 42854 124048 42938
rect 123728 42618 123770 42854
rect 124006 42618 124048 42854
rect 123728 42586 124048 42618
rect 154448 43174 154768 43206
rect 154448 42938 154490 43174
rect 154726 42938 154768 43174
rect 154448 42854 154768 42938
rect 154448 42618 154490 42854
rect 154726 42618 154768 42854
rect 154448 42586 154768 42618
rect 185168 43174 185488 43206
rect 185168 42938 185210 43174
rect 185446 42938 185488 43174
rect 185168 42854 185488 42938
rect 185168 42618 185210 42854
rect 185446 42618 185488 42854
rect 185168 42586 185488 42618
rect 215888 43174 216208 43206
rect 215888 42938 215930 43174
rect 216166 42938 216208 43174
rect 215888 42854 216208 42938
rect 215888 42618 215930 42854
rect 216166 42618 216208 42854
rect 215888 42586 216208 42618
rect 246608 43174 246928 43206
rect 246608 42938 246650 43174
rect 246886 42938 246928 43174
rect 246608 42854 246928 42938
rect 246608 42618 246650 42854
rect 246886 42618 246928 42854
rect 246608 42586 246928 42618
rect 277328 43174 277648 43206
rect 277328 42938 277370 43174
rect 277606 42938 277648 43174
rect 277328 42854 277648 42938
rect 277328 42618 277370 42854
rect 277606 42618 277648 42854
rect 277328 42586 277648 42618
rect 308048 43174 308368 43206
rect 308048 42938 308090 43174
rect 308326 42938 308368 43174
rect 308048 42854 308368 42938
rect 308048 42618 308090 42854
rect 308326 42618 308368 42854
rect 308048 42586 308368 42618
rect 338768 43174 339088 43206
rect 338768 42938 338810 43174
rect 339046 42938 339088 43174
rect 338768 42854 339088 42938
rect 338768 42618 338810 42854
rect 339046 42618 339088 42854
rect 338768 42586 339088 42618
rect 369488 43174 369808 43206
rect 369488 42938 369530 43174
rect 369766 42938 369808 43174
rect 369488 42854 369808 42938
rect 369488 42618 369530 42854
rect 369766 42618 369808 42854
rect 369488 42586 369808 42618
rect 400208 43174 400528 43206
rect 400208 42938 400250 43174
rect 400486 42938 400528 43174
rect 400208 42854 400528 42938
rect 400208 42618 400250 42854
rect 400486 42618 400528 42854
rect 400208 42586 400528 42618
rect 430928 43174 431248 43206
rect 430928 42938 430970 43174
rect 431206 42938 431248 43174
rect 430928 42854 431248 42938
rect 430928 42618 430970 42854
rect 431206 42618 431248 42854
rect 430928 42586 431248 42618
rect 461648 43174 461968 43206
rect 461648 42938 461690 43174
rect 461926 42938 461968 43174
rect 461648 42854 461968 42938
rect 461648 42618 461690 42854
rect 461926 42618 461968 42854
rect 461648 42586 461968 42618
rect 492368 43174 492688 43206
rect 492368 42938 492410 43174
rect 492646 42938 492688 43174
rect 492368 42854 492688 42938
rect 492368 42618 492410 42854
rect 492646 42618 492688 42854
rect 492368 42586 492688 42618
rect 523088 43174 523408 43206
rect 523088 42938 523130 43174
rect 523366 42938 523408 43174
rect 523088 42854 523408 42938
rect 523088 42618 523130 42854
rect 523366 42618 523408 42854
rect 523088 42586 523408 42618
rect 16208 39454 16528 39486
rect 16208 39218 16250 39454
rect 16486 39218 16528 39454
rect 16208 39134 16528 39218
rect 16208 38898 16250 39134
rect 16486 38898 16528 39134
rect 16208 38866 16528 38898
rect 46928 39454 47248 39486
rect 46928 39218 46970 39454
rect 47206 39218 47248 39454
rect 46928 39134 47248 39218
rect 46928 38898 46970 39134
rect 47206 38898 47248 39134
rect 46928 38866 47248 38898
rect 77648 39454 77968 39486
rect 77648 39218 77690 39454
rect 77926 39218 77968 39454
rect 77648 39134 77968 39218
rect 77648 38898 77690 39134
rect 77926 38898 77968 39134
rect 77648 38866 77968 38898
rect 108368 39454 108688 39486
rect 108368 39218 108410 39454
rect 108646 39218 108688 39454
rect 108368 39134 108688 39218
rect 108368 38898 108410 39134
rect 108646 38898 108688 39134
rect 108368 38866 108688 38898
rect 139088 39454 139408 39486
rect 139088 39218 139130 39454
rect 139366 39218 139408 39454
rect 139088 39134 139408 39218
rect 139088 38898 139130 39134
rect 139366 38898 139408 39134
rect 139088 38866 139408 38898
rect 169808 39454 170128 39486
rect 169808 39218 169850 39454
rect 170086 39218 170128 39454
rect 169808 39134 170128 39218
rect 169808 38898 169850 39134
rect 170086 38898 170128 39134
rect 169808 38866 170128 38898
rect 200528 39454 200848 39486
rect 200528 39218 200570 39454
rect 200806 39218 200848 39454
rect 200528 39134 200848 39218
rect 200528 38898 200570 39134
rect 200806 38898 200848 39134
rect 200528 38866 200848 38898
rect 231248 39454 231568 39486
rect 231248 39218 231290 39454
rect 231526 39218 231568 39454
rect 231248 39134 231568 39218
rect 231248 38898 231290 39134
rect 231526 38898 231568 39134
rect 231248 38866 231568 38898
rect 261968 39454 262288 39486
rect 261968 39218 262010 39454
rect 262246 39218 262288 39454
rect 261968 39134 262288 39218
rect 261968 38898 262010 39134
rect 262246 38898 262288 39134
rect 261968 38866 262288 38898
rect 292688 39454 293008 39486
rect 292688 39218 292730 39454
rect 292966 39218 293008 39454
rect 292688 39134 293008 39218
rect 292688 38898 292730 39134
rect 292966 38898 293008 39134
rect 292688 38866 293008 38898
rect 323408 39454 323728 39486
rect 323408 39218 323450 39454
rect 323686 39218 323728 39454
rect 323408 39134 323728 39218
rect 323408 38898 323450 39134
rect 323686 38898 323728 39134
rect 323408 38866 323728 38898
rect 354128 39454 354448 39486
rect 354128 39218 354170 39454
rect 354406 39218 354448 39454
rect 354128 39134 354448 39218
rect 354128 38898 354170 39134
rect 354406 38898 354448 39134
rect 354128 38866 354448 38898
rect 384848 39454 385168 39486
rect 384848 39218 384890 39454
rect 385126 39218 385168 39454
rect 384848 39134 385168 39218
rect 384848 38898 384890 39134
rect 385126 38898 385168 39134
rect 384848 38866 385168 38898
rect 415568 39454 415888 39486
rect 415568 39218 415610 39454
rect 415846 39218 415888 39454
rect 415568 39134 415888 39218
rect 415568 38898 415610 39134
rect 415846 38898 415888 39134
rect 415568 38866 415888 38898
rect 446288 39454 446608 39486
rect 446288 39218 446330 39454
rect 446566 39218 446608 39454
rect 446288 39134 446608 39218
rect 446288 38898 446330 39134
rect 446566 38898 446608 39134
rect 446288 38866 446608 38898
rect 477008 39454 477328 39486
rect 477008 39218 477050 39454
rect 477286 39218 477328 39454
rect 477008 39134 477328 39218
rect 477008 38898 477050 39134
rect 477286 38898 477328 39134
rect 477008 38866 477328 38898
rect 507728 39454 508048 39486
rect 507728 39218 507770 39454
rect 508006 39218 508048 39454
rect 507728 39134 508048 39218
rect 507728 38898 507770 39134
rect 508006 38898 508048 39134
rect 507728 38866 508048 38898
rect 538448 39454 538768 39486
rect 538448 39218 538490 39454
rect 538726 39218 538768 39454
rect 538448 39134 538768 39218
rect 538448 38898 538490 39134
rect 538726 38898 538768 39134
rect 538448 38866 538768 38898
rect 556674 18334 557294 53778
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 37794 3454 38414 13103
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 7174 42134 13103
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 10894 45854 13103
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 73794 3454 74414 13103
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 7174 78134 12068
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 10894 81854 13103
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 109794 3454 110414 13103
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 7174 114134 13103
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 10894 117854 13103
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 145794 3454 146414 13103
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 7174 150134 13103
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 10894 153854 13103
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 181794 3454 182414 13103
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 7174 186134 12068
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 10894 189854 13103
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 217794 3454 218414 13103
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 7174 222134 13103
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 10894 225854 13103
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 253794 3454 254414 13103
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 7174 258134 13103
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 10894 261854 13103
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 289794 3454 290414 13103
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 7174 294134 13103
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 10894 297854 13103
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 325794 3454 326414 13103
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 7174 330134 13103
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 10894 333854 13103
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 361794 3454 362414 13103
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 7174 366134 13103
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 10894 369854 12068
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 397794 3454 398414 13103
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 7174 402134 13103
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 10894 405854 13103
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 433794 3454 434414 13103
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 7174 438134 13103
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 10894 441854 13103
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 469794 3454 470414 13103
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 7174 474134 13103
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 10894 477854 12068
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 505794 3454 506414 13103
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 7174 510134 13103
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 10894 513854 13103
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 541794 3454 542414 13103
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 13103
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 10894 549854 13103
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 24146 710362 24382 710598
rect 24466 710362 24702 710598
rect 24146 710042 24382 710278
rect 24466 710042 24702 710278
rect 24146 673538 24382 673774
rect 24466 673538 24702 673774
rect 24146 673218 24382 673454
rect 24466 673218 24702 673454
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 52706 708442 52942 708678
rect 53026 708442 53262 708678
rect 52706 708122 52942 708358
rect 53026 708122 53262 708358
rect 52706 666098 52942 666334
rect 53026 666098 53262 666334
rect 52706 665778 52942 666014
rect 53026 665778 53262 666014
rect 56426 709402 56662 709638
rect 56746 709402 56982 709638
rect 56426 709082 56662 709318
rect 56746 709082 56982 709318
rect 56426 669818 56662 670054
rect 56746 669818 56982 670054
rect 56426 669498 56662 669734
rect 56746 669498 56982 669734
rect 60146 710362 60382 710598
rect 60466 710362 60702 710598
rect 60146 710042 60382 710278
rect 60466 710042 60702 710278
rect 60146 673538 60382 673774
rect 60466 673538 60702 673774
rect 60146 673218 60382 673454
rect 60466 673218 60702 673454
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 88706 708442 88942 708678
rect 89026 708442 89262 708678
rect 88706 708122 88942 708358
rect 89026 708122 89262 708358
rect 88706 666098 88942 666334
rect 89026 666098 89262 666334
rect 88706 665778 88942 666014
rect 89026 665778 89262 666014
rect 92426 709402 92662 709638
rect 92746 709402 92982 709638
rect 92426 709082 92662 709318
rect 92746 709082 92982 709318
rect 92426 669818 92662 670054
rect 92746 669818 92982 670054
rect 92426 669498 92662 669734
rect 92746 669498 92982 669734
rect 96146 710362 96382 710598
rect 96466 710362 96702 710598
rect 96146 710042 96382 710278
rect 96466 710042 96702 710278
rect 96146 673538 96382 673774
rect 96466 673538 96702 673774
rect 96146 673218 96382 673454
rect 96466 673218 96702 673454
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 124706 708442 124942 708678
rect 125026 708442 125262 708678
rect 124706 708122 124942 708358
rect 125026 708122 125262 708358
rect 124706 666098 124942 666334
rect 125026 666098 125262 666334
rect 124706 665778 124942 666014
rect 125026 665778 125262 666014
rect 128426 709402 128662 709638
rect 128746 709402 128982 709638
rect 128426 709082 128662 709318
rect 128746 709082 128982 709318
rect 128426 669818 128662 670054
rect 128746 669818 128982 670054
rect 128426 669498 128662 669734
rect 128746 669498 128982 669734
rect 132146 710362 132382 710598
rect 132466 710362 132702 710598
rect 132146 710042 132382 710278
rect 132466 710042 132702 710278
rect 132146 673538 132382 673774
rect 132466 673538 132702 673774
rect 132146 673218 132382 673454
rect 132466 673218 132702 673454
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 160706 708442 160942 708678
rect 161026 708442 161262 708678
rect 160706 708122 160942 708358
rect 161026 708122 161262 708358
rect 160706 666098 160942 666334
rect 161026 666098 161262 666334
rect 160706 665778 160942 666014
rect 161026 665778 161262 666014
rect 164426 709402 164662 709638
rect 164746 709402 164982 709638
rect 164426 709082 164662 709318
rect 164746 709082 164982 709318
rect 164426 669818 164662 670054
rect 164746 669818 164982 670054
rect 164426 669498 164662 669734
rect 164746 669498 164982 669734
rect 168146 710362 168382 710598
rect 168466 710362 168702 710598
rect 168146 710042 168382 710278
rect 168466 710042 168702 710278
rect 168146 673538 168382 673774
rect 168466 673538 168702 673774
rect 168146 673218 168382 673454
rect 168466 673218 168702 673454
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 196706 708442 196942 708678
rect 197026 708442 197262 708678
rect 196706 708122 196942 708358
rect 197026 708122 197262 708358
rect 196706 666098 196942 666334
rect 197026 666098 197262 666334
rect 196706 665778 196942 666014
rect 197026 665778 197262 666014
rect 200426 709402 200662 709638
rect 200746 709402 200982 709638
rect 200426 709082 200662 709318
rect 200746 709082 200982 709318
rect 200426 669818 200662 670054
rect 200746 669818 200982 670054
rect 200426 669498 200662 669734
rect 200746 669498 200982 669734
rect 204146 710362 204382 710598
rect 204466 710362 204702 710598
rect 204146 710042 204382 710278
rect 204466 710042 204702 710278
rect 204146 673538 204382 673774
rect 204466 673538 204702 673774
rect 204146 673218 204382 673454
rect 204466 673218 204702 673454
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 232706 708442 232942 708678
rect 233026 708442 233262 708678
rect 232706 708122 232942 708358
rect 233026 708122 233262 708358
rect 232706 666098 232942 666334
rect 233026 666098 233262 666334
rect 232706 665778 232942 666014
rect 233026 665778 233262 666014
rect 236426 709402 236662 709638
rect 236746 709402 236982 709638
rect 236426 709082 236662 709318
rect 236746 709082 236982 709318
rect 236426 669818 236662 670054
rect 236746 669818 236982 670054
rect 236426 669498 236662 669734
rect 236746 669498 236982 669734
rect 240146 710362 240382 710598
rect 240466 710362 240702 710598
rect 240146 710042 240382 710278
rect 240466 710042 240702 710278
rect 240146 673538 240382 673774
rect 240466 673538 240702 673774
rect 240146 673218 240382 673454
rect 240466 673218 240702 673454
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 268706 708442 268942 708678
rect 269026 708442 269262 708678
rect 268706 708122 268942 708358
rect 269026 708122 269262 708358
rect 268706 666098 268942 666334
rect 269026 666098 269262 666334
rect 268706 665778 268942 666014
rect 269026 665778 269262 666014
rect 272426 709402 272662 709638
rect 272746 709402 272982 709638
rect 272426 709082 272662 709318
rect 272746 709082 272982 709318
rect 272426 669818 272662 670054
rect 272746 669818 272982 670054
rect 272426 669498 272662 669734
rect 272746 669498 272982 669734
rect 276146 710362 276382 710598
rect 276466 710362 276702 710598
rect 276146 710042 276382 710278
rect 276466 710042 276702 710278
rect 276146 673538 276382 673774
rect 276466 673538 276702 673774
rect 276146 673218 276382 673454
rect 276466 673218 276702 673454
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 304706 708442 304942 708678
rect 305026 708442 305262 708678
rect 304706 708122 304942 708358
rect 305026 708122 305262 708358
rect 304706 666098 304942 666334
rect 305026 666098 305262 666334
rect 304706 665778 304942 666014
rect 305026 665778 305262 666014
rect 308426 709402 308662 709638
rect 308746 709402 308982 709638
rect 308426 709082 308662 709318
rect 308746 709082 308982 709318
rect 308426 669818 308662 670054
rect 308746 669818 308982 670054
rect 308426 669498 308662 669734
rect 308746 669498 308982 669734
rect 312146 710362 312382 710598
rect 312466 710362 312702 710598
rect 312146 710042 312382 710278
rect 312466 710042 312702 710278
rect 312146 673538 312382 673774
rect 312466 673538 312702 673774
rect 312146 673218 312382 673454
rect 312466 673218 312702 673454
rect 315866 711322 316102 711558
rect 316186 711322 316422 711558
rect 315866 711002 316102 711238
rect 316186 711002 316422 711238
rect 315866 677258 316102 677494
rect 316186 677258 316422 677494
rect 315866 676938 316102 677174
rect 316186 676938 316422 677174
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 340706 708442 340942 708678
rect 341026 708442 341262 708678
rect 340706 708122 340942 708358
rect 341026 708122 341262 708358
rect 340706 666098 340942 666334
rect 341026 666098 341262 666334
rect 340706 665778 340942 666014
rect 341026 665778 341262 666014
rect 344426 709402 344662 709638
rect 344746 709402 344982 709638
rect 344426 709082 344662 709318
rect 344746 709082 344982 709318
rect 344426 669818 344662 670054
rect 344746 669818 344982 670054
rect 344426 669498 344662 669734
rect 344746 669498 344982 669734
rect 348146 710362 348382 710598
rect 348466 710362 348702 710598
rect 348146 710042 348382 710278
rect 348466 710042 348702 710278
rect 348146 673538 348382 673774
rect 348466 673538 348702 673774
rect 348146 673218 348382 673454
rect 348466 673218 348702 673454
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 484706 708442 484942 708678
rect 485026 708442 485262 708678
rect 484706 708122 484942 708358
rect 485026 708122 485262 708358
rect 484706 666098 484942 666334
rect 485026 666098 485262 666334
rect 484706 665778 484942 666014
rect 485026 665778 485262 666014
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 31610 654938 31846 655174
rect 31610 654618 31846 654854
rect 62330 654938 62566 655174
rect 62330 654618 62566 654854
rect 93050 654938 93286 655174
rect 93050 654618 93286 654854
rect 123770 654938 124006 655174
rect 123770 654618 124006 654854
rect 154490 654938 154726 655174
rect 154490 654618 154726 654854
rect 185210 654938 185446 655174
rect 185210 654618 185446 654854
rect 215930 654938 216166 655174
rect 215930 654618 216166 654854
rect 246650 654938 246886 655174
rect 246650 654618 246886 654854
rect 277370 654938 277606 655174
rect 277370 654618 277606 654854
rect 308090 654938 308326 655174
rect 308090 654618 308326 654854
rect 338810 654938 339046 655174
rect 338810 654618 339046 654854
rect 369530 654938 369766 655174
rect 369530 654618 369766 654854
rect 400250 654938 400486 655174
rect 400250 654618 400486 654854
rect 430970 654938 431206 655174
rect 430970 654618 431206 654854
rect 461690 654938 461926 655174
rect 461690 654618 461926 654854
rect 492410 654938 492646 655174
rect 492410 654618 492646 654854
rect 523130 654938 523366 655174
rect 523130 654618 523366 654854
rect 16250 651218 16486 651454
rect 16250 650898 16486 651134
rect 46970 651218 47206 651454
rect 46970 650898 47206 651134
rect 77690 651218 77926 651454
rect 77690 650898 77926 651134
rect 108410 651218 108646 651454
rect 108410 650898 108646 651134
rect 139130 651218 139366 651454
rect 139130 650898 139366 651134
rect 169850 651218 170086 651454
rect 169850 650898 170086 651134
rect 200570 651218 200806 651454
rect 200570 650898 200806 651134
rect 231290 651218 231526 651454
rect 231290 650898 231526 651134
rect 262010 651218 262246 651454
rect 262010 650898 262246 651134
rect 292730 651218 292966 651454
rect 292730 650898 292966 651134
rect 323450 651218 323686 651454
rect 323450 650898 323686 651134
rect 354170 651218 354406 651454
rect 354170 650898 354406 651134
rect 384890 651218 385126 651454
rect 384890 650898 385126 651134
rect 415610 651218 415846 651454
rect 415610 650898 415846 651134
rect 446330 651218 446566 651454
rect 446330 650898 446566 651134
rect 477050 651218 477286 651454
rect 477050 650898 477286 651134
rect 507770 651218 508006 651454
rect 507770 650898 508006 651134
rect 538490 651218 538726 651454
rect 538490 650898 538726 651134
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 31610 618938 31846 619174
rect 31610 618618 31846 618854
rect 62330 618938 62566 619174
rect 62330 618618 62566 618854
rect 93050 618938 93286 619174
rect 93050 618618 93286 618854
rect 123770 618938 124006 619174
rect 123770 618618 124006 618854
rect 154490 618938 154726 619174
rect 154490 618618 154726 618854
rect 185210 618938 185446 619174
rect 185210 618618 185446 618854
rect 215930 618938 216166 619174
rect 215930 618618 216166 618854
rect 246650 618938 246886 619174
rect 246650 618618 246886 618854
rect 277370 618938 277606 619174
rect 277370 618618 277606 618854
rect 308090 618938 308326 619174
rect 308090 618618 308326 618854
rect 338810 618938 339046 619174
rect 338810 618618 339046 618854
rect 369530 618938 369766 619174
rect 369530 618618 369766 618854
rect 400250 618938 400486 619174
rect 400250 618618 400486 618854
rect 430970 618938 431206 619174
rect 430970 618618 431206 618854
rect 461690 618938 461926 619174
rect 461690 618618 461926 618854
rect 492410 618938 492646 619174
rect 492410 618618 492646 618854
rect 523130 618938 523366 619174
rect 523130 618618 523366 618854
rect 16250 615218 16486 615454
rect 16250 614898 16486 615134
rect 46970 615218 47206 615454
rect 46970 614898 47206 615134
rect 77690 615218 77926 615454
rect 77690 614898 77926 615134
rect 108410 615218 108646 615454
rect 108410 614898 108646 615134
rect 139130 615218 139366 615454
rect 139130 614898 139366 615134
rect 169850 615218 170086 615454
rect 169850 614898 170086 615134
rect 200570 615218 200806 615454
rect 200570 614898 200806 615134
rect 231290 615218 231526 615454
rect 231290 614898 231526 615134
rect 262010 615218 262246 615454
rect 262010 614898 262246 615134
rect 292730 615218 292966 615454
rect 292730 614898 292966 615134
rect 323450 615218 323686 615454
rect 323450 614898 323686 615134
rect 354170 615218 354406 615454
rect 354170 614898 354406 615134
rect 384890 615218 385126 615454
rect 384890 614898 385126 615134
rect 415610 615218 415846 615454
rect 415610 614898 415846 615134
rect 446330 615218 446566 615454
rect 446330 614898 446566 615134
rect 477050 615218 477286 615454
rect 477050 614898 477286 615134
rect 507770 615218 508006 615454
rect 507770 614898 508006 615134
rect 538490 615218 538726 615454
rect 538490 614898 538726 615134
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 31610 582938 31846 583174
rect 31610 582618 31846 582854
rect 62330 582938 62566 583174
rect 62330 582618 62566 582854
rect 93050 582938 93286 583174
rect 93050 582618 93286 582854
rect 123770 582938 124006 583174
rect 123770 582618 124006 582854
rect 154490 582938 154726 583174
rect 154490 582618 154726 582854
rect 185210 582938 185446 583174
rect 185210 582618 185446 582854
rect 215930 582938 216166 583174
rect 215930 582618 216166 582854
rect 246650 582938 246886 583174
rect 246650 582618 246886 582854
rect 277370 582938 277606 583174
rect 277370 582618 277606 582854
rect 308090 582938 308326 583174
rect 308090 582618 308326 582854
rect 338810 582938 339046 583174
rect 338810 582618 339046 582854
rect 369530 582938 369766 583174
rect 369530 582618 369766 582854
rect 400250 582938 400486 583174
rect 400250 582618 400486 582854
rect 430970 582938 431206 583174
rect 430970 582618 431206 582854
rect 461690 582938 461926 583174
rect 461690 582618 461926 582854
rect 492410 582938 492646 583174
rect 492410 582618 492646 582854
rect 523130 582938 523366 583174
rect 523130 582618 523366 582854
rect 16250 579218 16486 579454
rect 16250 578898 16486 579134
rect 46970 579218 47206 579454
rect 46970 578898 47206 579134
rect 77690 579218 77926 579454
rect 77690 578898 77926 579134
rect 108410 579218 108646 579454
rect 108410 578898 108646 579134
rect 139130 579218 139366 579454
rect 139130 578898 139366 579134
rect 169850 579218 170086 579454
rect 169850 578898 170086 579134
rect 200570 579218 200806 579454
rect 200570 578898 200806 579134
rect 231290 579218 231526 579454
rect 231290 578898 231526 579134
rect 262010 579218 262246 579454
rect 262010 578898 262246 579134
rect 292730 579218 292966 579454
rect 292730 578898 292966 579134
rect 323450 579218 323686 579454
rect 323450 578898 323686 579134
rect 354170 579218 354406 579454
rect 354170 578898 354406 579134
rect 384890 579218 385126 579454
rect 384890 578898 385126 579134
rect 415610 579218 415846 579454
rect 415610 578898 415846 579134
rect 446330 579218 446566 579454
rect 446330 578898 446566 579134
rect 477050 579218 477286 579454
rect 477050 578898 477286 579134
rect 507770 579218 508006 579454
rect 507770 578898 508006 579134
rect 538490 579218 538726 579454
rect 538490 578898 538726 579134
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 31610 546938 31846 547174
rect 31610 546618 31846 546854
rect 62330 546938 62566 547174
rect 62330 546618 62566 546854
rect 93050 546938 93286 547174
rect 93050 546618 93286 546854
rect 123770 546938 124006 547174
rect 123770 546618 124006 546854
rect 154490 546938 154726 547174
rect 154490 546618 154726 546854
rect 185210 546938 185446 547174
rect 185210 546618 185446 546854
rect 215930 546938 216166 547174
rect 215930 546618 216166 546854
rect 246650 546938 246886 547174
rect 246650 546618 246886 546854
rect 277370 546938 277606 547174
rect 277370 546618 277606 546854
rect 308090 546938 308326 547174
rect 308090 546618 308326 546854
rect 338810 546938 339046 547174
rect 338810 546618 339046 546854
rect 369530 546938 369766 547174
rect 369530 546618 369766 546854
rect 400250 546938 400486 547174
rect 400250 546618 400486 546854
rect 430970 546938 431206 547174
rect 430970 546618 431206 546854
rect 461690 546938 461926 547174
rect 461690 546618 461926 546854
rect 492410 546938 492646 547174
rect 492410 546618 492646 546854
rect 523130 546938 523366 547174
rect 523130 546618 523366 546854
rect 16250 543218 16486 543454
rect 16250 542898 16486 543134
rect 46970 543218 47206 543454
rect 46970 542898 47206 543134
rect 77690 543218 77926 543454
rect 77690 542898 77926 543134
rect 108410 543218 108646 543454
rect 108410 542898 108646 543134
rect 139130 543218 139366 543454
rect 139130 542898 139366 543134
rect 169850 543218 170086 543454
rect 169850 542898 170086 543134
rect 200570 543218 200806 543454
rect 200570 542898 200806 543134
rect 231290 543218 231526 543454
rect 231290 542898 231526 543134
rect 262010 543218 262246 543454
rect 262010 542898 262246 543134
rect 292730 543218 292966 543454
rect 292730 542898 292966 543134
rect 323450 543218 323686 543454
rect 323450 542898 323686 543134
rect 354170 543218 354406 543454
rect 354170 542898 354406 543134
rect 384890 543218 385126 543454
rect 384890 542898 385126 543134
rect 415610 543218 415846 543454
rect 415610 542898 415846 543134
rect 446330 543218 446566 543454
rect 446330 542898 446566 543134
rect 477050 543218 477286 543454
rect 477050 542898 477286 543134
rect 507770 543218 508006 543454
rect 507770 542898 508006 543134
rect 538490 543218 538726 543454
rect 538490 542898 538726 543134
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 31610 510938 31846 511174
rect 31610 510618 31846 510854
rect 62330 510938 62566 511174
rect 62330 510618 62566 510854
rect 93050 510938 93286 511174
rect 93050 510618 93286 510854
rect 123770 510938 124006 511174
rect 123770 510618 124006 510854
rect 154490 510938 154726 511174
rect 154490 510618 154726 510854
rect 185210 510938 185446 511174
rect 185210 510618 185446 510854
rect 215930 510938 216166 511174
rect 215930 510618 216166 510854
rect 246650 510938 246886 511174
rect 246650 510618 246886 510854
rect 277370 510938 277606 511174
rect 277370 510618 277606 510854
rect 308090 510938 308326 511174
rect 308090 510618 308326 510854
rect 338810 510938 339046 511174
rect 338810 510618 339046 510854
rect 369530 510938 369766 511174
rect 369530 510618 369766 510854
rect 400250 510938 400486 511174
rect 400250 510618 400486 510854
rect 430970 510938 431206 511174
rect 430970 510618 431206 510854
rect 461690 510938 461926 511174
rect 461690 510618 461926 510854
rect 492410 510938 492646 511174
rect 492410 510618 492646 510854
rect 523130 510938 523366 511174
rect 523130 510618 523366 510854
rect 16250 507218 16486 507454
rect 16250 506898 16486 507134
rect 46970 507218 47206 507454
rect 46970 506898 47206 507134
rect 77690 507218 77926 507454
rect 77690 506898 77926 507134
rect 108410 507218 108646 507454
rect 108410 506898 108646 507134
rect 139130 507218 139366 507454
rect 139130 506898 139366 507134
rect 169850 507218 170086 507454
rect 169850 506898 170086 507134
rect 200570 507218 200806 507454
rect 200570 506898 200806 507134
rect 231290 507218 231526 507454
rect 231290 506898 231526 507134
rect 262010 507218 262246 507454
rect 262010 506898 262246 507134
rect 292730 507218 292966 507454
rect 292730 506898 292966 507134
rect 323450 507218 323686 507454
rect 323450 506898 323686 507134
rect 354170 507218 354406 507454
rect 354170 506898 354406 507134
rect 384890 507218 385126 507454
rect 384890 506898 385126 507134
rect 415610 507218 415846 507454
rect 415610 506898 415846 507134
rect 446330 507218 446566 507454
rect 446330 506898 446566 507134
rect 477050 507218 477286 507454
rect 477050 506898 477286 507134
rect 507770 507218 508006 507454
rect 507770 506898 508006 507134
rect 538490 507218 538726 507454
rect 538490 506898 538726 507134
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 31610 474938 31846 475174
rect 31610 474618 31846 474854
rect 62330 474938 62566 475174
rect 62330 474618 62566 474854
rect 93050 474938 93286 475174
rect 93050 474618 93286 474854
rect 123770 474938 124006 475174
rect 123770 474618 124006 474854
rect 154490 474938 154726 475174
rect 154490 474618 154726 474854
rect 185210 474938 185446 475174
rect 185210 474618 185446 474854
rect 215930 474938 216166 475174
rect 215930 474618 216166 474854
rect 246650 474938 246886 475174
rect 246650 474618 246886 474854
rect 277370 474938 277606 475174
rect 277370 474618 277606 474854
rect 308090 474938 308326 475174
rect 308090 474618 308326 474854
rect 338810 474938 339046 475174
rect 338810 474618 339046 474854
rect 369530 474938 369766 475174
rect 369530 474618 369766 474854
rect 400250 474938 400486 475174
rect 400250 474618 400486 474854
rect 430970 474938 431206 475174
rect 430970 474618 431206 474854
rect 461690 474938 461926 475174
rect 461690 474618 461926 474854
rect 492410 474938 492646 475174
rect 492410 474618 492646 474854
rect 523130 474938 523366 475174
rect 523130 474618 523366 474854
rect 16250 471218 16486 471454
rect 16250 470898 16486 471134
rect 46970 471218 47206 471454
rect 46970 470898 47206 471134
rect 77690 471218 77926 471454
rect 77690 470898 77926 471134
rect 108410 471218 108646 471454
rect 108410 470898 108646 471134
rect 139130 471218 139366 471454
rect 139130 470898 139366 471134
rect 169850 471218 170086 471454
rect 169850 470898 170086 471134
rect 200570 471218 200806 471454
rect 200570 470898 200806 471134
rect 231290 471218 231526 471454
rect 231290 470898 231526 471134
rect 262010 471218 262246 471454
rect 262010 470898 262246 471134
rect 292730 471218 292966 471454
rect 292730 470898 292966 471134
rect 323450 471218 323686 471454
rect 323450 470898 323686 471134
rect 354170 471218 354406 471454
rect 354170 470898 354406 471134
rect 384890 471218 385126 471454
rect 384890 470898 385126 471134
rect 415610 471218 415846 471454
rect 415610 470898 415846 471134
rect 446330 471218 446566 471454
rect 446330 470898 446566 471134
rect 477050 471218 477286 471454
rect 477050 470898 477286 471134
rect 507770 471218 508006 471454
rect 507770 470898 508006 471134
rect 538490 471218 538726 471454
rect 538490 470898 538726 471134
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 31610 438938 31846 439174
rect 31610 438618 31846 438854
rect 62330 438938 62566 439174
rect 62330 438618 62566 438854
rect 93050 438938 93286 439174
rect 93050 438618 93286 438854
rect 123770 438938 124006 439174
rect 123770 438618 124006 438854
rect 154490 438938 154726 439174
rect 154490 438618 154726 438854
rect 185210 438938 185446 439174
rect 185210 438618 185446 438854
rect 215930 438938 216166 439174
rect 215930 438618 216166 438854
rect 246650 438938 246886 439174
rect 246650 438618 246886 438854
rect 277370 438938 277606 439174
rect 277370 438618 277606 438854
rect 308090 438938 308326 439174
rect 308090 438618 308326 438854
rect 338810 438938 339046 439174
rect 338810 438618 339046 438854
rect 369530 438938 369766 439174
rect 369530 438618 369766 438854
rect 400250 438938 400486 439174
rect 400250 438618 400486 438854
rect 430970 438938 431206 439174
rect 430970 438618 431206 438854
rect 461690 438938 461926 439174
rect 461690 438618 461926 438854
rect 492410 438938 492646 439174
rect 492410 438618 492646 438854
rect 523130 438938 523366 439174
rect 523130 438618 523366 438854
rect 16250 435218 16486 435454
rect 16250 434898 16486 435134
rect 46970 435218 47206 435454
rect 46970 434898 47206 435134
rect 77690 435218 77926 435454
rect 77690 434898 77926 435134
rect 108410 435218 108646 435454
rect 108410 434898 108646 435134
rect 139130 435218 139366 435454
rect 139130 434898 139366 435134
rect 169850 435218 170086 435454
rect 169850 434898 170086 435134
rect 200570 435218 200806 435454
rect 200570 434898 200806 435134
rect 231290 435218 231526 435454
rect 231290 434898 231526 435134
rect 262010 435218 262246 435454
rect 262010 434898 262246 435134
rect 292730 435218 292966 435454
rect 292730 434898 292966 435134
rect 323450 435218 323686 435454
rect 323450 434898 323686 435134
rect 354170 435218 354406 435454
rect 354170 434898 354406 435134
rect 384890 435218 385126 435454
rect 384890 434898 385126 435134
rect 415610 435218 415846 435454
rect 415610 434898 415846 435134
rect 446330 435218 446566 435454
rect 446330 434898 446566 435134
rect 477050 435218 477286 435454
rect 477050 434898 477286 435134
rect 507770 435218 508006 435454
rect 507770 434898 508006 435134
rect 538490 435218 538726 435454
rect 538490 434898 538726 435134
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 31610 402938 31846 403174
rect 31610 402618 31846 402854
rect 62330 402938 62566 403174
rect 62330 402618 62566 402854
rect 93050 402938 93286 403174
rect 93050 402618 93286 402854
rect 123770 402938 124006 403174
rect 123770 402618 124006 402854
rect 154490 402938 154726 403174
rect 154490 402618 154726 402854
rect 185210 402938 185446 403174
rect 185210 402618 185446 402854
rect 215930 402938 216166 403174
rect 215930 402618 216166 402854
rect 246650 402938 246886 403174
rect 246650 402618 246886 402854
rect 277370 402938 277606 403174
rect 277370 402618 277606 402854
rect 308090 402938 308326 403174
rect 308090 402618 308326 402854
rect 338810 402938 339046 403174
rect 338810 402618 339046 402854
rect 369530 402938 369766 403174
rect 369530 402618 369766 402854
rect 400250 402938 400486 403174
rect 400250 402618 400486 402854
rect 430970 402938 431206 403174
rect 430970 402618 431206 402854
rect 461690 402938 461926 403174
rect 461690 402618 461926 402854
rect 492410 402938 492646 403174
rect 492410 402618 492646 402854
rect 523130 402938 523366 403174
rect 523130 402618 523366 402854
rect 16250 399218 16486 399454
rect 16250 398898 16486 399134
rect 46970 399218 47206 399454
rect 46970 398898 47206 399134
rect 77690 399218 77926 399454
rect 77690 398898 77926 399134
rect 108410 399218 108646 399454
rect 108410 398898 108646 399134
rect 139130 399218 139366 399454
rect 139130 398898 139366 399134
rect 169850 399218 170086 399454
rect 169850 398898 170086 399134
rect 200570 399218 200806 399454
rect 200570 398898 200806 399134
rect 231290 399218 231526 399454
rect 231290 398898 231526 399134
rect 262010 399218 262246 399454
rect 262010 398898 262246 399134
rect 292730 399218 292966 399454
rect 292730 398898 292966 399134
rect 323450 399218 323686 399454
rect 323450 398898 323686 399134
rect 354170 399218 354406 399454
rect 354170 398898 354406 399134
rect 384890 399218 385126 399454
rect 384890 398898 385126 399134
rect 415610 399218 415846 399454
rect 415610 398898 415846 399134
rect 446330 399218 446566 399454
rect 446330 398898 446566 399134
rect 477050 399218 477286 399454
rect 477050 398898 477286 399134
rect 507770 399218 508006 399454
rect 507770 398898 508006 399134
rect 538490 399218 538726 399454
rect 538490 398898 538726 399134
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 556706 378098 556942 378334
rect 557026 378098 557262 378334
rect 556706 377778 556942 378014
rect 557026 377778 557262 378014
rect 31610 366938 31846 367174
rect 31610 366618 31846 366854
rect 62330 366938 62566 367174
rect 62330 366618 62566 366854
rect 93050 366938 93286 367174
rect 93050 366618 93286 366854
rect 123770 366938 124006 367174
rect 123770 366618 124006 366854
rect 154490 366938 154726 367174
rect 154490 366618 154726 366854
rect 185210 366938 185446 367174
rect 185210 366618 185446 366854
rect 215930 366938 216166 367174
rect 215930 366618 216166 366854
rect 246650 366938 246886 367174
rect 246650 366618 246886 366854
rect 277370 366938 277606 367174
rect 277370 366618 277606 366854
rect 308090 366938 308326 367174
rect 308090 366618 308326 366854
rect 338810 366938 339046 367174
rect 338810 366618 339046 366854
rect 369530 366938 369766 367174
rect 369530 366618 369766 366854
rect 400250 366938 400486 367174
rect 400250 366618 400486 366854
rect 430970 366938 431206 367174
rect 430970 366618 431206 366854
rect 461690 366938 461926 367174
rect 461690 366618 461926 366854
rect 492410 366938 492646 367174
rect 492410 366618 492646 366854
rect 523130 366938 523366 367174
rect 523130 366618 523366 366854
rect 16250 363218 16486 363454
rect 16250 362898 16486 363134
rect 46970 363218 47206 363454
rect 46970 362898 47206 363134
rect 77690 363218 77926 363454
rect 77690 362898 77926 363134
rect 108410 363218 108646 363454
rect 108410 362898 108646 363134
rect 139130 363218 139366 363454
rect 139130 362898 139366 363134
rect 169850 363218 170086 363454
rect 169850 362898 170086 363134
rect 200570 363218 200806 363454
rect 200570 362898 200806 363134
rect 231290 363218 231526 363454
rect 231290 362898 231526 363134
rect 262010 363218 262246 363454
rect 262010 362898 262246 363134
rect 292730 363218 292966 363454
rect 292730 362898 292966 363134
rect 323450 363218 323686 363454
rect 323450 362898 323686 363134
rect 354170 363218 354406 363454
rect 354170 362898 354406 363134
rect 384890 363218 385126 363454
rect 384890 362898 385126 363134
rect 415610 363218 415846 363454
rect 415610 362898 415846 363134
rect 446330 363218 446566 363454
rect 446330 362898 446566 363134
rect 477050 363218 477286 363454
rect 477050 362898 477286 363134
rect 507770 363218 508006 363454
rect 507770 362898 508006 363134
rect 538490 363218 538726 363454
rect 538490 362898 538726 363134
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 31610 330938 31846 331174
rect 31610 330618 31846 330854
rect 62330 330938 62566 331174
rect 62330 330618 62566 330854
rect 93050 330938 93286 331174
rect 93050 330618 93286 330854
rect 123770 330938 124006 331174
rect 123770 330618 124006 330854
rect 154490 330938 154726 331174
rect 154490 330618 154726 330854
rect 185210 330938 185446 331174
rect 185210 330618 185446 330854
rect 215930 330938 216166 331174
rect 215930 330618 216166 330854
rect 246650 330938 246886 331174
rect 246650 330618 246886 330854
rect 277370 330938 277606 331174
rect 277370 330618 277606 330854
rect 308090 330938 308326 331174
rect 308090 330618 308326 330854
rect 338810 330938 339046 331174
rect 338810 330618 339046 330854
rect 369530 330938 369766 331174
rect 369530 330618 369766 330854
rect 400250 330938 400486 331174
rect 400250 330618 400486 330854
rect 430970 330938 431206 331174
rect 430970 330618 431206 330854
rect 461690 330938 461926 331174
rect 461690 330618 461926 330854
rect 492410 330938 492646 331174
rect 492410 330618 492646 330854
rect 523130 330938 523366 331174
rect 523130 330618 523366 330854
rect 16250 327218 16486 327454
rect 16250 326898 16486 327134
rect 46970 327218 47206 327454
rect 46970 326898 47206 327134
rect 77690 327218 77926 327454
rect 77690 326898 77926 327134
rect 108410 327218 108646 327454
rect 108410 326898 108646 327134
rect 139130 327218 139366 327454
rect 139130 326898 139366 327134
rect 169850 327218 170086 327454
rect 169850 326898 170086 327134
rect 200570 327218 200806 327454
rect 200570 326898 200806 327134
rect 231290 327218 231526 327454
rect 231290 326898 231526 327134
rect 262010 327218 262246 327454
rect 262010 326898 262246 327134
rect 292730 327218 292966 327454
rect 292730 326898 292966 327134
rect 323450 327218 323686 327454
rect 323450 326898 323686 327134
rect 354170 327218 354406 327454
rect 354170 326898 354406 327134
rect 384890 327218 385126 327454
rect 384890 326898 385126 327134
rect 415610 327218 415846 327454
rect 415610 326898 415846 327134
rect 446330 327218 446566 327454
rect 446330 326898 446566 327134
rect 477050 327218 477286 327454
rect 477050 326898 477286 327134
rect 507770 327218 508006 327454
rect 507770 326898 508006 327134
rect 538490 327218 538726 327454
rect 538490 326898 538726 327134
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 31610 294938 31846 295174
rect 31610 294618 31846 294854
rect 62330 294938 62566 295174
rect 62330 294618 62566 294854
rect 93050 294938 93286 295174
rect 93050 294618 93286 294854
rect 123770 294938 124006 295174
rect 123770 294618 124006 294854
rect 154490 294938 154726 295174
rect 154490 294618 154726 294854
rect 185210 294938 185446 295174
rect 185210 294618 185446 294854
rect 215930 294938 216166 295174
rect 215930 294618 216166 294854
rect 246650 294938 246886 295174
rect 246650 294618 246886 294854
rect 277370 294938 277606 295174
rect 277370 294618 277606 294854
rect 308090 294938 308326 295174
rect 308090 294618 308326 294854
rect 338810 294938 339046 295174
rect 338810 294618 339046 294854
rect 369530 294938 369766 295174
rect 369530 294618 369766 294854
rect 400250 294938 400486 295174
rect 400250 294618 400486 294854
rect 430970 294938 431206 295174
rect 430970 294618 431206 294854
rect 461690 294938 461926 295174
rect 461690 294618 461926 294854
rect 492410 294938 492646 295174
rect 492410 294618 492646 294854
rect 523130 294938 523366 295174
rect 523130 294618 523366 294854
rect 16250 291218 16486 291454
rect 16250 290898 16486 291134
rect 46970 291218 47206 291454
rect 46970 290898 47206 291134
rect 77690 291218 77926 291454
rect 77690 290898 77926 291134
rect 108410 291218 108646 291454
rect 108410 290898 108646 291134
rect 139130 291218 139366 291454
rect 139130 290898 139366 291134
rect 169850 291218 170086 291454
rect 169850 290898 170086 291134
rect 200570 291218 200806 291454
rect 200570 290898 200806 291134
rect 231290 291218 231526 291454
rect 231290 290898 231526 291134
rect 262010 291218 262246 291454
rect 262010 290898 262246 291134
rect 292730 291218 292966 291454
rect 292730 290898 292966 291134
rect 323450 291218 323686 291454
rect 323450 290898 323686 291134
rect 354170 291218 354406 291454
rect 354170 290898 354406 291134
rect 384890 291218 385126 291454
rect 384890 290898 385126 291134
rect 415610 291218 415846 291454
rect 415610 290898 415846 291134
rect 446330 291218 446566 291454
rect 446330 290898 446566 291134
rect 477050 291218 477286 291454
rect 477050 290898 477286 291134
rect 507770 291218 508006 291454
rect 507770 290898 508006 291134
rect 538490 291218 538726 291454
rect 538490 290898 538726 291134
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 31610 258938 31846 259174
rect 31610 258618 31846 258854
rect 62330 258938 62566 259174
rect 62330 258618 62566 258854
rect 93050 258938 93286 259174
rect 93050 258618 93286 258854
rect 123770 258938 124006 259174
rect 123770 258618 124006 258854
rect 154490 258938 154726 259174
rect 154490 258618 154726 258854
rect 185210 258938 185446 259174
rect 185210 258618 185446 258854
rect 215930 258938 216166 259174
rect 215930 258618 216166 258854
rect 246650 258938 246886 259174
rect 246650 258618 246886 258854
rect 277370 258938 277606 259174
rect 277370 258618 277606 258854
rect 308090 258938 308326 259174
rect 308090 258618 308326 258854
rect 338810 258938 339046 259174
rect 338810 258618 339046 258854
rect 369530 258938 369766 259174
rect 369530 258618 369766 258854
rect 400250 258938 400486 259174
rect 400250 258618 400486 258854
rect 430970 258938 431206 259174
rect 430970 258618 431206 258854
rect 461690 258938 461926 259174
rect 461690 258618 461926 258854
rect 492410 258938 492646 259174
rect 492410 258618 492646 258854
rect 523130 258938 523366 259174
rect 523130 258618 523366 258854
rect 16250 255218 16486 255454
rect 16250 254898 16486 255134
rect 46970 255218 47206 255454
rect 46970 254898 47206 255134
rect 77690 255218 77926 255454
rect 77690 254898 77926 255134
rect 108410 255218 108646 255454
rect 108410 254898 108646 255134
rect 139130 255218 139366 255454
rect 139130 254898 139366 255134
rect 169850 255218 170086 255454
rect 169850 254898 170086 255134
rect 200570 255218 200806 255454
rect 200570 254898 200806 255134
rect 231290 255218 231526 255454
rect 231290 254898 231526 255134
rect 262010 255218 262246 255454
rect 262010 254898 262246 255134
rect 292730 255218 292966 255454
rect 292730 254898 292966 255134
rect 323450 255218 323686 255454
rect 323450 254898 323686 255134
rect 354170 255218 354406 255454
rect 354170 254898 354406 255134
rect 384890 255218 385126 255454
rect 384890 254898 385126 255134
rect 415610 255218 415846 255454
rect 415610 254898 415846 255134
rect 446330 255218 446566 255454
rect 446330 254898 446566 255134
rect 477050 255218 477286 255454
rect 477050 254898 477286 255134
rect 507770 255218 508006 255454
rect 507770 254898 508006 255134
rect 538490 255218 538726 255454
rect 538490 254898 538726 255134
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 31610 222938 31846 223174
rect 31610 222618 31846 222854
rect 62330 222938 62566 223174
rect 62330 222618 62566 222854
rect 93050 222938 93286 223174
rect 93050 222618 93286 222854
rect 123770 222938 124006 223174
rect 123770 222618 124006 222854
rect 154490 222938 154726 223174
rect 154490 222618 154726 222854
rect 185210 222938 185446 223174
rect 185210 222618 185446 222854
rect 215930 222938 216166 223174
rect 215930 222618 216166 222854
rect 246650 222938 246886 223174
rect 246650 222618 246886 222854
rect 277370 222938 277606 223174
rect 277370 222618 277606 222854
rect 308090 222938 308326 223174
rect 308090 222618 308326 222854
rect 338810 222938 339046 223174
rect 338810 222618 339046 222854
rect 369530 222938 369766 223174
rect 369530 222618 369766 222854
rect 400250 222938 400486 223174
rect 400250 222618 400486 222854
rect 430970 222938 431206 223174
rect 430970 222618 431206 222854
rect 461690 222938 461926 223174
rect 461690 222618 461926 222854
rect 492410 222938 492646 223174
rect 492410 222618 492646 222854
rect 523130 222938 523366 223174
rect 523130 222618 523366 222854
rect 16250 219218 16486 219454
rect 16250 218898 16486 219134
rect 46970 219218 47206 219454
rect 46970 218898 47206 219134
rect 77690 219218 77926 219454
rect 77690 218898 77926 219134
rect 108410 219218 108646 219454
rect 108410 218898 108646 219134
rect 139130 219218 139366 219454
rect 139130 218898 139366 219134
rect 169850 219218 170086 219454
rect 169850 218898 170086 219134
rect 200570 219218 200806 219454
rect 200570 218898 200806 219134
rect 231290 219218 231526 219454
rect 231290 218898 231526 219134
rect 262010 219218 262246 219454
rect 262010 218898 262246 219134
rect 292730 219218 292966 219454
rect 292730 218898 292966 219134
rect 323450 219218 323686 219454
rect 323450 218898 323686 219134
rect 354170 219218 354406 219454
rect 354170 218898 354406 219134
rect 384890 219218 385126 219454
rect 384890 218898 385126 219134
rect 415610 219218 415846 219454
rect 415610 218898 415846 219134
rect 446330 219218 446566 219454
rect 446330 218898 446566 219134
rect 477050 219218 477286 219454
rect 477050 218898 477286 219134
rect 507770 219218 508006 219454
rect 507770 218898 508006 219134
rect 538490 219218 538726 219454
rect 538490 218898 538726 219134
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 31610 186938 31846 187174
rect 31610 186618 31846 186854
rect 62330 186938 62566 187174
rect 62330 186618 62566 186854
rect 93050 186938 93286 187174
rect 93050 186618 93286 186854
rect 123770 186938 124006 187174
rect 123770 186618 124006 186854
rect 154490 186938 154726 187174
rect 154490 186618 154726 186854
rect 185210 186938 185446 187174
rect 185210 186618 185446 186854
rect 215930 186938 216166 187174
rect 215930 186618 216166 186854
rect 246650 186938 246886 187174
rect 246650 186618 246886 186854
rect 277370 186938 277606 187174
rect 277370 186618 277606 186854
rect 308090 186938 308326 187174
rect 308090 186618 308326 186854
rect 338810 186938 339046 187174
rect 338810 186618 339046 186854
rect 369530 186938 369766 187174
rect 369530 186618 369766 186854
rect 400250 186938 400486 187174
rect 400250 186618 400486 186854
rect 430970 186938 431206 187174
rect 430970 186618 431206 186854
rect 461690 186938 461926 187174
rect 461690 186618 461926 186854
rect 492410 186938 492646 187174
rect 492410 186618 492646 186854
rect 523130 186938 523366 187174
rect 523130 186618 523366 186854
rect 16250 183218 16486 183454
rect 16250 182898 16486 183134
rect 46970 183218 47206 183454
rect 46970 182898 47206 183134
rect 77690 183218 77926 183454
rect 77690 182898 77926 183134
rect 108410 183218 108646 183454
rect 108410 182898 108646 183134
rect 139130 183218 139366 183454
rect 139130 182898 139366 183134
rect 169850 183218 170086 183454
rect 169850 182898 170086 183134
rect 200570 183218 200806 183454
rect 200570 182898 200806 183134
rect 231290 183218 231526 183454
rect 231290 182898 231526 183134
rect 262010 183218 262246 183454
rect 262010 182898 262246 183134
rect 292730 183218 292966 183454
rect 292730 182898 292966 183134
rect 323450 183218 323686 183454
rect 323450 182898 323686 183134
rect 354170 183218 354406 183454
rect 354170 182898 354406 183134
rect 384890 183218 385126 183454
rect 384890 182898 385126 183134
rect 415610 183218 415846 183454
rect 415610 182898 415846 183134
rect 446330 183218 446566 183454
rect 446330 182898 446566 183134
rect 477050 183218 477286 183454
rect 477050 182898 477286 183134
rect 507770 183218 508006 183454
rect 507770 182898 508006 183134
rect 538490 183218 538726 183454
rect 538490 182898 538726 183134
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 31610 150938 31846 151174
rect 31610 150618 31846 150854
rect 62330 150938 62566 151174
rect 62330 150618 62566 150854
rect 93050 150938 93286 151174
rect 93050 150618 93286 150854
rect 123770 150938 124006 151174
rect 123770 150618 124006 150854
rect 154490 150938 154726 151174
rect 154490 150618 154726 150854
rect 185210 150938 185446 151174
rect 185210 150618 185446 150854
rect 215930 150938 216166 151174
rect 215930 150618 216166 150854
rect 246650 150938 246886 151174
rect 246650 150618 246886 150854
rect 277370 150938 277606 151174
rect 277370 150618 277606 150854
rect 308090 150938 308326 151174
rect 308090 150618 308326 150854
rect 338810 150938 339046 151174
rect 338810 150618 339046 150854
rect 369530 150938 369766 151174
rect 369530 150618 369766 150854
rect 400250 150938 400486 151174
rect 400250 150618 400486 150854
rect 430970 150938 431206 151174
rect 430970 150618 431206 150854
rect 461690 150938 461926 151174
rect 461690 150618 461926 150854
rect 492410 150938 492646 151174
rect 492410 150618 492646 150854
rect 523130 150938 523366 151174
rect 523130 150618 523366 150854
rect 16250 147218 16486 147454
rect 16250 146898 16486 147134
rect 46970 147218 47206 147454
rect 46970 146898 47206 147134
rect 77690 147218 77926 147454
rect 77690 146898 77926 147134
rect 108410 147218 108646 147454
rect 108410 146898 108646 147134
rect 139130 147218 139366 147454
rect 139130 146898 139366 147134
rect 169850 147218 170086 147454
rect 169850 146898 170086 147134
rect 200570 147218 200806 147454
rect 200570 146898 200806 147134
rect 231290 147218 231526 147454
rect 231290 146898 231526 147134
rect 262010 147218 262246 147454
rect 262010 146898 262246 147134
rect 292730 147218 292966 147454
rect 292730 146898 292966 147134
rect 323450 147218 323686 147454
rect 323450 146898 323686 147134
rect 354170 147218 354406 147454
rect 354170 146898 354406 147134
rect 384890 147218 385126 147454
rect 384890 146898 385126 147134
rect 415610 147218 415846 147454
rect 415610 146898 415846 147134
rect 446330 147218 446566 147454
rect 446330 146898 446566 147134
rect 477050 147218 477286 147454
rect 477050 146898 477286 147134
rect 507770 147218 508006 147454
rect 507770 146898 508006 147134
rect 538490 147218 538726 147454
rect 538490 146898 538726 147134
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 31610 114938 31846 115174
rect 31610 114618 31846 114854
rect 62330 114938 62566 115174
rect 62330 114618 62566 114854
rect 93050 114938 93286 115174
rect 93050 114618 93286 114854
rect 123770 114938 124006 115174
rect 123770 114618 124006 114854
rect 154490 114938 154726 115174
rect 154490 114618 154726 114854
rect 185210 114938 185446 115174
rect 185210 114618 185446 114854
rect 215930 114938 216166 115174
rect 215930 114618 216166 114854
rect 246650 114938 246886 115174
rect 246650 114618 246886 114854
rect 277370 114938 277606 115174
rect 277370 114618 277606 114854
rect 308090 114938 308326 115174
rect 308090 114618 308326 114854
rect 338810 114938 339046 115174
rect 338810 114618 339046 114854
rect 369530 114938 369766 115174
rect 369530 114618 369766 114854
rect 400250 114938 400486 115174
rect 400250 114618 400486 114854
rect 430970 114938 431206 115174
rect 430970 114618 431206 114854
rect 461690 114938 461926 115174
rect 461690 114618 461926 114854
rect 492410 114938 492646 115174
rect 492410 114618 492646 114854
rect 523130 114938 523366 115174
rect 523130 114618 523366 114854
rect 16250 111218 16486 111454
rect 16250 110898 16486 111134
rect 46970 111218 47206 111454
rect 46970 110898 47206 111134
rect 77690 111218 77926 111454
rect 77690 110898 77926 111134
rect 108410 111218 108646 111454
rect 108410 110898 108646 111134
rect 139130 111218 139366 111454
rect 139130 110898 139366 111134
rect 169850 111218 170086 111454
rect 169850 110898 170086 111134
rect 200570 111218 200806 111454
rect 200570 110898 200806 111134
rect 231290 111218 231526 111454
rect 231290 110898 231526 111134
rect 262010 111218 262246 111454
rect 262010 110898 262246 111134
rect 292730 111218 292966 111454
rect 292730 110898 292966 111134
rect 323450 111218 323686 111454
rect 323450 110898 323686 111134
rect 354170 111218 354406 111454
rect 354170 110898 354406 111134
rect 384890 111218 385126 111454
rect 384890 110898 385126 111134
rect 415610 111218 415846 111454
rect 415610 110898 415846 111134
rect 446330 111218 446566 111454
rect 446330 110898 446566 111134
rect 477050 111218 477286 111454
rect 477050 110898 477286 111134
rect 507770 111218 508006 111454
rect 507770 110898 508006 111134
rect 538490 111218 538726 111454
rect 538490 110898 538726 111134
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 31610 78938 31846 79174
rect 31610 78618 31846 78854
rect 62330 78938 62566 79174
rect 62330 78618 62566 78854
rect 93050 78938 93286 79174
rect 93050 78618 93286 78854
rect 123770 78938 124006 79174
rect 123770 78618 124006 78854
rect 154490 78938 154726 79174
rect 154490 78618 154726 78854
rect 185210 78938 185446 79174
rect 185210 78618 185446 78854
rect 215930 78938 216166 79174
rect 215930 78618 216166 78854
rect 246650 78938 246886 79174
rect 246650 78618 246886 78854
rect 277370 78938 277606 79174
rect 277370 78618 277606 78854
rect 308090 78938 308326 79174
rect 308090 78618 308326 78854
rect 338810 78938 339046 79174
rect 338810 78618 339046 78854
rect 369530 78938 369766 79174
rect 369530 78618 369766 78854
rect 400250 78938 400486 79174
rect 400250 78618 400486 78854
rect 430970 78938 431206 79174
rect 430970 78618 431206 78854
rect 461690 78938 461926 79174
rect 461690 78618 461926 78854
rect 492410 78938 492646 79174
rect 492410 78618 492646 78854
rect 523130 78938 523366 79174
rect 523130 78618 523366 78854
rect 16250 75218 16486 75454
rect 16250 74898 16486 75134
rect 46970 75218 47206 75454
rect 46970 74898 47206 75134
rect 77690 75218 77926 75454
rect 77690 74898 77926 75134
rect 108410 75218 108646 75454
rect 108410 74898 108646 75134
rect 139130 75218 139366 75454
rect 139130 74898 139366 75134
rect 169850 75218 170086 75454
rect 169850 74898 170086 75134
rect 200570 75218 200806 75454
rect 200570 74898 200806 75134
rect 231290 75218 231526 75454
rect 231290 74898 231526 75134
rect 262010 75218 262246 75454
rect 262010 74898 262246 75134
rect 292730 75218 292966 75454
rect 292730 74898 292966 75134
rect 323450 75218 323686 75454
rect 323450 74898 323686 75134
rect 354170 75218 354406 75454
rect 354170 74898 354406 75134
rect 384890 75218 385126 75454
rect 384890 74898 385126 75134
rect 415610 75218 415846 75454
rect 415610 74898 415846 75134
rect 446330 75218 446566 75454
rect 446330 74898 446566 75134
rect 477050 75218 477286 75454
rect 477050 74898 477286 75134
rect 507770 75218 508006 75454
rect 507770 74898 508006 75134
rect 538490 75218 538726 75454
rect 538490 74898 538726 75134
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 31610 42938 31846 43174
rect 31610 42618 31846 42854
rect 62330 42938 62566 43174
rect 62330 42618 62566 42854
rect 93050 42938 93286 43174
rect 93050 42618 93286 42854
rect 123770 42938 124006 43174
rect 123770 42618 124006 42854
rect 154490 42938 154726 43174
rect 154490 42618 154726 42854
rect 185210 42938 185446 43174
rect 185210 42618 185446 42854
rect 215930 42938 216166 43174
rect 215930 42618 216166 42854
rect 246650 42938 246886 43174
rect 246650 42618 246886 42854
rect 277370 42938 277606 43174
rect 277370 42618 277606 42854
rect 308090 42938 308326 43174
rect 308090 42618 308326 42854
rect 338810 42938 339046 43174
rect 338810 42618 339046 42854
rect 369530 42938 369766 43174
rect 369530 42618 369766 42854
rect 400250 42938 400486 43174
rect 400250 42618 400486 42854
rect 430970 42938 431206 43174
rect 430970 42618 431206 42854
rect 461690 42938 461926 43174
rect 461690 42618 461926 42854
rect 492410 42938 492646 43174
rect 492410 42618 492646 42854
rect 523130 42938 523366 43174
rect 523130 42618 523366 42854
rect 16250 39218 16486 39454
rect 16250 38898 16486 39134
rect 46970 39218 47206 39454
rect 46970 38898 47206 39134
rect 77690 39218 77926 39454
rect 77690 38898 77926 39134
rect 108410 39218 108646 39454
rect 108410 38898 108646 39134
rect 139130 39218 139366 39454
rect 139130 38898 139366 39134
rect 169850 39218 170086 39454
rect 169850 38898 170086 39134
rect 200570 39218 200806 39454
rect 200570 38898 200806 39134
rect 231290 39218 231526 39454
rect 231290 38898 231526 39134
rect 262010 39218 262246 39454
rect 262010 38898 262246 39134
rect 292730 39218 292966 39454
rect 292730 38898 292966 39134
rect 323450 39218 323686 39454
rect 323450 38898 323686 39134
rect 354170 39218 354406 39454
rect 354170 38898 354406 39134
rect 384890 39218 385126 39454
rect 384890 38898 385126 39134
rect 415610 39218 415846 39454
rect 415610 38898 415846 39134
rect 446330 39218 446566 39454
rect 446330 38898 446566 39134
rect 477050 39218 477286 39454
rect 477050 38898 477286 39134
rect 507770 39218 508006 39454
rect 507770 38898 508006 39134
rect 538490 39218 538726 39454
rect 538490 38898 538726 39134
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 31610 655174
rect 31846 654938 62330 655174
rect 62566 654938 93050 655174
rect 93286 654938 123770 655174
rect 124006 654938 154490 655174
rect 154726 654938 185210 655174
rect 185446 654938 215930 655174
rect 216166 654938 246650 655174
rect 246886 654938 277370 655174
rect 277606 654938 308090 655174
rect 308326 654938 338810 655174
rect 339046 654938 369530 655174
rect 369766 654938 400250 655174
rect 400486 654938 430970 655174
rect 431206 654938 461690 655174
rect 461926 654938 492410 655174
rect 492646 654938 523130 655174
rect 523366 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 31610 654854
rect 31846 654618 62330 654854
rect 62566 654618 93050 654854
rect 93286 654618 123770 654854
rect 124006 654618 154490 654854
rect 154726 654618 185210 654854
rect 185446 654618 215930 654854
rect 216166 654618 246650 654854
rect 246886 654618 277370 654854
rect 277606 654618 308090 654854
rect 308326 654618 338810 654854
rect 339046 654618 369530 654854
rect 369766 654618 400250 654854
rect 400486 654618 430970 654854
rect 431206 654618 461690 654854
rect 461926 654618 492410 654854
rect 492646 654618 523130 654854
rect 523366 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 16250 651454
rect 16486 651218 46970 651454
rect 47206 651218 77690 651454
rect 77926 651218 108410 651454
rect 108646 651218 139130 651454
rect 139366 651218 169850 651454
rect 170086 651218 200570 651454
rect 200806 651218 231290 651454
rect 231526 651218 262010 651454
rect 262246 651218 292730 651454
rect 292966 651218 323450 651454
rect 323686 651218 354170 651454
rect 354406 651218 384890 651454
rect 385126 651218 415610 651454
rect 415846 651218 446330 651454
rect 446566 651218 477050 651454
rect 477286 651218 507770 651454
rect 508006 651218 538490 651454
rect 538726 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 16250 651134
rect 16486 650898 46970 651134
rect 47206 650898 77690 651134
rect 77926 650898 108410 651134
rect 108646 650898 139130 651134
rect 139366 650898 169850 651134
rect 170086 650898 200570 651134
rect 200806 650898 231290 651134
rect 231526 650898 262010 651134
rect 262246 650898 292730 651134
rect 292966 650898 323450 651134
rect 323686 650898 354170 651134
rect 354406 650898 384890 651134
rect 385126 650898 415610 651134
rect 415846 650898 446330 651134
rect 446566 650898 477050 651134
rect 477286 650898 507770 651134
rect 508006 650898 538490 651134
rect 538726 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 31610 619174
rect 31846 618938 62330 619174
rect 62566 618938 93050 619174
rect 93286 618938 123770 619174
rect 124006 618938 154490 619174
rect 154726 618938 185210 619174
rect 185446 618938 215930 619174
rect 216166 618938 246650 619174
rect 246886 618938 277370 619174
rect 277606 618938 308090 619174
rect 308326 618938 338810 619174
rect 339046 618938 369530 619174
rect 369766 618938 400250 619174
rect 400486 618938 430970 619174
rect 431206 618938 461690 619174
rect 461926 618938 492410 619174
rect 492646 618938 523130 619174
rect 523366 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 31610 618854
rect 31846 618618 62330 618854
rect 62566 618618 93050 618854
rect 93286 618618 123770 618854
rect 124006 618618 154490 618854
rect 154726 618618 185210 618854
rect 185446 618618 215930 618854
rect 216166 618618 246650 618854
rect 246886 618618 277370 618854
rect 277606 618618 308090 618854
rect 308326 618618 338810 618854
rect 339046 618618 369530 618854
rect 369766 618618 400250 618854
rect 400486 618618 430970 618854
rect 431206 618618 461690 618854
rect 461926 618618 492410 618854
rect 492646 618618 523130 618854
rect 523366 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 16250 615454
rect 16486 615218 46970 615454
rect 47206 615218 77690 615454
rect 77926 615218 108410 615454
rect 108646 615218 139130 615454
rect 139366 615218 169850 615454
rect 170086 615218 200570 615454
rect 200806 615218 231290 615454
rect 231526 615218 262010 615454
rect 262246 615218 292730 615454
rect 292966 615218 323450 615454
rect 323686 615218 354170 615454
rect 354406 615218 384890 615454
rect 385126 615218 415610 615454
rect 415846 615218 446330 615454
rect 446566 615218 477050 615454
rect 477286 615218 507770 615454
rect 508006 615218 538490 615454
rect 538726 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 16250 615134
rect 16486 614898 46970 615134
rect 47206 614898 77690 615134
rect 77926 614898 108410 615134
rect 108646 614898 139130 615134
rect 139366 614898 169850 615134
rect 170086 614898 200570 615134
rect 200806 614898 231290 615134
rect 231526 614898 262010 615134
rect 262246 614898 292730 615134
rect 292966 614898 323450 615134
rect 323686 614898 354170 615134
rect 354406 614898 384890 615134
rect 385126 614898 415610 615134
rect 415846 614898 446330 615134
rect 446566 614898 477050 615134
rect 477286 614898 507770 615134
rect 508006 614898 538490 615134
rect 538726 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 31610 583174
rect 31846 582938 62330 583174
rect 62566 582938 93050 583174
rect 93286 582938 123770 583174
rect 124006 582938 154490 583174
rect 154726 582938 185210 583174
rect 185446 582938 215930 583174
rect 216166 582938 246650 583174
rect 246886 582938 277370 583174
rect 277606 582938 308090 583174
rect 308326 582938 338810 583174
rect 339046 582938 369530 583174
rect 369766 582938 400250 583174
rect 400486 582938 430970 583174
rect 431206 582938 461690 583174
rect 461926 582938 492410 583174
rect 492646 582938 523130 583174
rect 523366 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 31610 582854
rect 31846 582618 62330 582854
rect 62566 582618 93050 582854
rect 93286 582618 123770 582854
rect 124006 582618 154490 582854
rect 154726 582618 185210 582854
rect 185446 582618 215930 582854
rect 216166 582618 246650 582854
rect 246886 582618 277370 582854
rect 277606 582618 308090 582854
rect 308326 582618 338810 582854
rect 339046 582618 369530 582854
rect 369766 582618 400250 582854
rect 400486 582618 430970 582854
rect 431206 582618 461690 582854
rect 461926 582618 492410 582854
rect 492646 582618 523130 582854
rect 523366 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 16250 579454
rect 16486 579218 46970 579454
rect 47206 579218 77690 579454
rect 77926 579218 108410 579454
rect 108646 579218 139130 579454
rect 139366 579218 169850 579454
rect 170086 579218 200570 579454
rect 200806 579218 231290 579454
rect 231526 579218 262010 579454
rect 262246 579218 292730 579454
rect 292966 579218 323450 579454
rect 323686 579218 354170 579454
rect 354406 579218 384890 579454
rect 385126 579218 415610 579454
rect 415846 579218 446330 579454
rect 446566 579218 477050 579454
rect 477286 579218 507770 579454
rect 508006 579218 538490 579454
rect 538726 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 16250 579134
rect 16486 578898 46970 579134
rect 47206 578898 77690 579134
rect 77926 578898 108410 579134
rect 108646 578898 139130 579134
rect 139366 578898 169850 579134
rect 170086 578898 200570 579134
rect 200806 578898 231290 579134
rect 231526 578898 262010 579134
rect 262246 578898 292730 579134
rect 292966 578898 323450 579134
rect 323686 578898 354170 579134
rect 354406 578898 384890 579134
rect 385126 578898 415610 579134
rect 415846 578898 446330 579134
rect 446566 578898 477050 579134
rect 477286 578898 507770 579134
rect 508006 578898 538490 579134
rect 538726 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 31610 547174
rect 31846 546938 62330 547174
rect 62566 546938 93050 547174
rect 93286 546938 123770 547174
rect 124006 546938 154490 547174
rect 154726 546938 185210 547174
rect 185446 546938 215930 547174
rect 216166 546938 246650 547174
rect 246886 546938 277370 547174
rect 277606 546938 308090 547174
rect 308326 546938 338810 547174
rect 339046 546938 369530 547174
rect 369766 546938 400250 547174
rect 400486 546938 430970 547174
rect 431206 546938 461690 547174
rect 461926 546938 492410 547174
rect 492646 546938 523130 547174
rect 523366 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 31610 546854
rect 31846 546618 62330 546854
rect 62566 546618 93050 546854
rect 93286 546618 123770 546854
rect 124006 546618 154490 546854
rect 154726 546618 185210 546854
rect 185446 546618 215930 546854
rect 216166 546618 246650 546854
rect 246886 546618 277370 546854
rect 277606 546618 308090 546854
rect 308326 546618 338810 546854
rect 339046 546618 369530 546854
rect 369766 546618 400250 546854
rect 400486 546618 430970 546854
rect 431206 546618 461690 546854
rect 461926 546618 492410 546854
rect 492646 546618 523130 546854
rect 523366 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 16250 543454
rect 16486 543218 46970 543454
rect 47206 543218 77690 543454
rect 77926 543218 108410 543454
rect 108646 543218 139130 543454
rect 139366 543218 169850 543454
rect 170086 543218 200570 543454
rect 200806 543218 231290 543454
rect 231526 543218 262010 543454
rect 262246 543218 292730 543454
rect 292966 543218 323450 543454
rect 323686 543218 354170 543454
rect 354406 543218 384890 543454
rect 385126 543218 415610 543454
rect 415846 543218 446330 543454
rect 446566 543218 477050 543454
rect 477286 543218 507770 543454
rect 508006 543218 538490 543454
rect 538726 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 16250 543134
rect 16486 542898 46970 543134
rect 47206 542898 77690 543134
rect 77926 542898 108410 543134
rect 108646 542898 139130 543134
rect 139366 542898 169850 543134
rect 170086 542898 200570 543134
rect 200806 542898 231290 543134
rect 231526 542898 262010 543134
rect 262246 542898 292730 543134
rect 292966 542898 323450 543134
rect 323686 542898 354170 543134
rect 354406 542898 384890 543134
rect 385126 542898 415610 543134
rect 415846 542898 446330 543134
rect 446566 542898 477050 543134
rect 477286 542898 507770 543134
rect 508006 542898 538490 543134
rect 538726 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 31610 511174
rect 31846 510938 62330 511174
rect 62566 510938 93050 511174
rect 93286 510938 123770 511174
rect 124006 510938 154490 511174
rect 154726 510938 185210 511174
rect 185446 510938 215930 511174
rect 216166 510938 246650 511174
rect 246886 510938 277370 511174
rect 277606 510938 308090 511174
rect 308326 510938 338810 511174
rect 339046 510938 369530 511174
rect 369766 510938 400250 511174
rect 400486 510938 430970 511174
rect 431206 510938 461690 511174
rect 461926 510938 492410 511174
rect 492646 510938 523130 511174
rect 523366 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 31610 510854
rect 31846 510618 62330 510854
rect 62566 510618 93050 510854
rect 93286 510618 123770 510854
rect 124006 510618 154490 510854
rect 154726 510618 185210 510854
rect 185446 510618 215930 510854
rect 216166 510618 246650 510854
rect 246886 510618 277370 510854
rect 277606 510618 308090 510854
rect 308326 510618 338810 510854
rect 339046 510618 369530 510854
rect 369766 510618 400250 510854
rect 400486 510618 430970 510854
rect 431206 510618 461690 510854
rect 461926 510618 492410 510854
rect 492646 510618 523130 510854
rect 523366 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 16250 507454
rect 16486 507218 46970 507454
rect 47206 507218 77690 507454
rect 77926 507218 108410 507454
rect 108646 507218 139130 507454
rect 139366 507218 169850 507454
rect 170086 507218 200570 507454
rect 200806 507218 231290 507454
rect 231526 507218 262010 507454
rect 262246 507218 292730 507454
rect 292966 507218 323450 507454
rect 323686 507218 354170 507454
rect 354406 507218 384890 507454
rect 385126 507218 415610 507454
rect 415846 507218 446330 507454
rect 446566 507218 477050 507454
rect 477286 507218 507770 507454
rect 508006 507218 538490 507454
rect 538726 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 16250 507134
rect 16486 506898 46970 507134
rect 47206 506898 77690 507134
rect 77926 506898 108410 507134
rect 108646 506898 139130 507134
rect 139366 506898 169850 507134
rect 170086 506898 200570 507134
rect 200806 506898 231290 507134
rect 231526 506898 262010 507134
rect 262246 506898 292730 507134
rect 292966 506898 323450 507134
rect 323686 506898 354170 507134
rect 354406 506898 384890 507134
rect 385126 506898 415610 507134
rect 415846 506898 446330 507134
rect 446566 506898 477050 507134
rect 477286 506898 507770 507134
rect 508006 506898 538490 507134
rect 538726 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 31610 475174
rect 31846 474938 62330 475174
rect 62566 474938 93050 475174
rect 93286 474938 123770 475174
rect 124006 474938 154490 475174
rect 154726 474938 185210 475174
rect 185446 474938 215930 475174
rect 216166 474938 246650 475174
rect 246886 474938 277370 475174
rect 277606 474938 308090 475174
rect 308326 474938 338810 475174
rect 339046 474938 369530 475174
rect 369766 474938 400250 475174
rect 400486 474938 430970 475174
rect 431206 474938 461690 475174
rect 461926 474938 492410 475174
rect 492646 474938 523130 475174
rect 523366 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 31610 474854
rect 31846 474618 62330 474854
rect 62566 474618 93050 474854
rect 93286 474618 123770 474854
rect 124006 474618 154490 474854
rect 154726 474618 185210 474854
rect 185446 474618 215930 474854
rect 216166 474618 246650 474854
rect 246886 474618 277370 474854
rect 277606 474618 308090 474854
rect 308326 474618 338810 474854
rect 339046 474618 369530 474854
rect 369766 474618 400250 474854
rect 400486 474618 430970 474854
rect 431206 474618 461690 474854
rect 461926 474618 492410 474854
rect 492646 474618 523130 474854
rect 523366 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 16250 471454
rect 16486 471218 46970 471454
rect 47206 471218 77690 471454
rect 77926 471218 108410 471454
rect 108646 471218 139130 471454
rect 139366 471218 169850 471454
rect 170086 471218 200570 471454
rect 200806 471218 231290 471454
rect 231526 471218 262010 471454
rect 262246 471218 292730 471454
rect 292966 471218 323450 471454
rect 323686 471218 354170 471454
rect 354406 471218 384890 471454
rect 385126 471218 415610 471454
rect 415846 471218 446330 471454
rect 446566 471218 477050 471454
rect 477286 471218 507770 471454
rect 508006 471218 538490 471454
rect 538726 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 16250 471134
rect 16486 470898 46970 471134
rect 47206 470898 77690 471134
rect 77926 470898 108410 471134
rect 108646 470898 139130 471134
rect 139366 470898 169850 471134
rect 170086 470898 200570 471134
rect 200806 470898 231290 471134
rect 231526 470898 262010 471134
rect 262246 470898 292730 471134
rect 292966 470898 323450 471134
rect 323686 470898 354170 471134
rect 354406 470898 384890 471134
rect 385126 470898 415610 471134
rect 415846 470898 446330 471134
rect 446566 470898 477050 471134
rect 477286 470898 507770 471134
rect 508006 470898 538490 471134
rect 538726 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 31610 439174
rect 31846 438938 62330 439174
rect 62566 438938 93050 439174
rect 93286 438938 123770 439174
rect 124006 438938 154490 439174
rect 154726 438938 185210 439174
rect 185446 438938 215930 439174
rect 216166 438938 246650 439174
rect 246886 438938 277370 439174
rect 277606 438938 308090 439174
rect 308326 438938 338810 439174
rect 339046 438938 369530 439174
rect 369766 438938 400250 439174
rect 400486 438938 430970 439174
rect 431206 438938 461690 439174
rect 461926 438938 492410 439174
rect 492646 438938 523130 439174
rect 523366 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 31610 438854
rect 31846 438618 62330 438854
rect 62566 438618 93050 438854
rect 93286 438618 123770 438854
rect 124006 438618 154490 438854
rect 154726 438618 185210 438854
rect 185446 438618 215930 438854
rect 216166 438618 246650 438854
rect 246886 438618 277370 438854
rect 277606 438618 308090 438854
rect 308326 438618 338810 438854
rect 339046 438618 369530 438854
rect 369766 438618 400250 438854
rect 400486 438618 430970 438854
rect 431206 438618 461690 438854
rect 461926 438618 492410 438854
rect 492646 438618 523130 438854
rect 523366 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 16250 435454
rect 16486 435218 46970 435454
rect 47206 435218 77690 435454
rect 77926 435218 108410 435454
rect 108646 435218 139130 435454
rect 139366 435218 169850 435454
rect 170086 435218 200570 435454
rect 200806 435218 231290 435454
rect 231526 435218 262010 435454
rect 262246 435218 292730 435454
rect 292966 435218 323450 435454
rect 323686 435218 354170 435454
rect 354406 435218 384890 435454
rect 385126 435218 415610 435454
rect 415846 435218 446330 435454
rect 446566 435218 477050 435454
rect 477286 435218 507770 435454
rect 508006 435218 538490 435454
rect 538726 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 16250 435134
rect 16486 434898 46970 435134
rect 47206 434898 77690 435134
rect 77926 434898 108410 435134
rect 108646 434898 139130 435134
rect 139366 434898 169850 435134
rect 170086 434898 200570 435134
rect 200806 434898 231290 435134
rect 231526 434898 262010 435134
rect 262246 434898 292730 435134
rect 292966 434898 323450 435134
rect 323686 434898 354170 435134
rect 354406 434898 384890 435134
rect 385126 434898 415610 435134
rect 415846 434898 446330 435134
rect 446566 434898 477050 435134
rect 477286 434898 507770 435134
rect 508006 434898 538490 435134
rect 538726 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 31610 403174
rect 31846 402938 62330 403174
rect 62566 402938 93050 403174
rect 93286 402938 123770 403174
rect 124006 402938 154490 403174
rect 154726 402938 185210 403174
rect 185446 402938 215930 403174
rect 216166 402938 246650 403174
rect 246886 402938 277370 403174
rect 277606 402938 308090 403174
rect 308326 402938 338810 403174
rect 339046 402938 369530 403174
rect 369766 402938 400250 403174
rect 400486 402938 430970 403174
rect 431206 402938 461690 403174
rect 461926 402938 492410 403174
rect 492646 402938 523130 403174
rect 523366 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 31610 402854
rect 31846 402618 62330 402854
rect 62566 402618 93050 402854
rect 93286 402618 123770 402854
rect 124006 402618 154490 402854
rect 154726 402618 185210 402854
rect 185446 402618 215930 402854
rect 216166 402618 246650 402854
rect 246886 402618 277370 402854
rect 277606 402618 308090 402854
rect 308326 402618 338810 402854
rect 339046 402618 369530 402854
rect 369766 402618 400250 402854
rect 400486 402618 430970 402854
rect 431206 402618 461690 402854
rect 461926 402618 492410 402854
rect 492646 402618 523130 402854
rect 523366 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 16250 399454
rect 16486 399218 46970 399454
rect 47206 399218 77690 399454
rect 77926 399218 108410 399454
rect 108646 399218 139130 399454
rect 139366 399218 169850 399454
rect 170086 399218 200570 399454
rect 200806 399218 231290 399454
rect 231526 399218 262010 399454
rect 262246 399218 292730 399454
rect 292966 399218 323450 399454
rect 323686 399218 354170 399454
rect 354406 399218 384890 399454
rect 385126 399218 415610 399454
rect 415846 399218 446330 399454
rect 446566 399218 477050 399454
rect 477286 399218 507770 399454
rect 508006 399218 538490 399454
rect 538726 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 16250 399134
rect 16486 398898 46970 399134
rect 47206 398898 77690 399134
rect 77926 398898 108410 399134
rect 108646 398898 139130 399134
rect 139366 398898 169850 399134
rect 170086 398898 200570 399134
rect 200806 398898 231290 399134
rect 231526 398898 262010 399134
rect 262246 398898 292730 399134
rect 292966 398898 323450 399134
rect 323686 398898 354170 399134
rect 354406 398898 384890 399134
rect 385126 398898 415610 399134
rect 415846 398898 446330 399134
rect 446566 398898 477050 399134
rect 477286 398898 507770 399134
rect 508006 398898 538490 399134
rect 538726 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 31610 367174
rect 31846 366938 62330 367174
rect 62566 366938 93050 367174
rect 93286 366938 123770 367174
rect 124006 366938 154490 367174
rect 154726 366938 185210 367174
rect 185446 366938 215930 367174
rect 216166 366938 246650 367174
rect 246886 366938 277370 367174
rect 277606 366938 308090 367174
rect 308326 366938 338810 367174
rect 339046 366938 369530 367174
rect 369766 366938 400250 367174
rect 400486 366938 430970 367174
rect 431206 366938 461690 367174
rect 461926 366938 492410 367174
rect 492646 366938 523130 367174
rect 523366 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 31610 366854
rect 31846 366618 62330 366854
rect 62566 366618 93050 366854
rect 93286 366618 123770 366854
rect 124006 366618 154490 366854
rect 154726 366618 185210 366854
rect 185446 366618 215930 366854
rect 216166 366618 246650 366854
rect 246886 366618 277370 366854
rect 277606 366618 308090 366854
rect 308326 366618 338810 366854
rect 339046 366618 369530 366854
rect 369766 366618 400250 366854
rect 400486 366618 430970 366854
rect 431206 366618 461690 366854
rect 461926 366618 492410 366854
rect 492646 366618 523130 366854
rect 523366 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 16250 363454
rect 16486 363218 46970 363454
rect 47206 363218 77690 363454
rect 77926 363218 108410 363454
rect 108646 363218 139130 363454
rect 139366 363218 169850 363454
rect 170086 363218 200570 363454
rect 200806 363218 231290 363454
rect 231526 363218 262010 363454
rect 262246 363218 292730 363454
rect 292966 363218 323450 363454
rect 323686 363218 354170 363454
rect 354406 363218 384890 363454
rect 385126 363218 415610 363454
rect 415846 363218 446330 363454
rect 446566 363218 477050 363454
rect 477286 363218 507770 363454
rect 508006 363218 538490 363454
rect 538726 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 16250 363134
rect 16486 362898 46970 363134
rect 47206 362898 77690 363134
rect 77926 362898 108410 363134
rect 108646 362898 139130 363134
rect 139366 362898 169850 363134
rect 170086 362898 200570 363134
rect 200806 362898 231290 363134
rect 231526 362898 262010 363134
rect 262246 362898 292730 363134
rect 292966 362898 323450 363134
rect 323686 362898 354170 363134
rect 354406 362898 384890 363134
rect 385126 362898 415610 363134
rect 415846 362898 446330 363134
rect 446566 362898 477050 363134
rect 477286 362898 507770 363134
rect 508006 362898 538490 363134
rect 538726 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 31610 331174
rect 31846 330938 62330 331174
rect 62566 330938 93050 331174
rect 93286 330938 123770 331174
rect 124006 330938 154490 331174
rect 154726 330938 185210 331174
rect 185446 330938 215930 331174
rect 216166 330938 246650 331174
rect 246886 330938 277370 331174
rect 277606 330938 308090 331174
rect 308326 330938 338810 331174
rect 339046 330938 369530 331174
rect 369766 330938 400250 331174
rect 400486 330938 430970 331174
rect 431206 330938 461690 331174
rect 461926 330938 492410 331174
rect 492646 330938 523130 331174
rect 523366 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 31610 330854
rect 31846 330618 62330 330854
rect 62566 330618 93050 330854
rect 93286 330618 123770 330854
rect 124006 330618 154490 330854
rect 154726 330618 185210 330854
rect 185446 330618 215930 330854
rect 216166 330618 246650 330854
rect 246886 330618 277370 330854
rect 277606 330618 308090 330854
rect 308326 330618 338810 330854
rect 339046 330618 369530 330854
rect 369766 330618 400250 330854
rect 400486 330618 430970 330854
rect 431206 330618 461690 330854
rect 461926 330618 492410 330854
rect 492646 330618 523130 330854
rect 523366 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 16250 327454
rect 16486 327218 46970 327454
rect 47206 327218 77690 327454
rect 77926 327218 108410 327454
rect 108646 327218 139130 327454
rect 139366 327218 169850 327454
rect 170086 327218 200570 327454
rect 200806 327218 231290 327454
rect 231526 327218 262010 327454
rect 262246 327218 292730 327454
rect 292966 327218 323450 327454
rect 323686 327218 354170 327454
rect 354406 327218 384890 327454
rect 385126 327218 415610 327454
rect 415846 327218 446330 327454
rect 446566 327218 477050 327454
rect 477286 327218 507770 327454
rect 508006 327218 538490 327454
rect 538726 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 16250 327134
rect 16486 326898 46970 327134
rect 47206 326898 77690 327134
rect 77926 326898 108410 327134
rect 108646 326898 139130 327134
rect 139366 326898 169850 327134
rect 170086 326898 200570 327134
rect 200806 326898 231290 327134
rect 231526 326898 262010 327134
rect 262246 326898 292730 327134
rect 292966 326898 323450 327134
rect 323686 326898 354170 327134
rect 354406 326898 384890 327134
rect 385126 326898 415610 327134
rect 415846 326898 446330 327134
rect 446566 326898 477050 327134
rect 477286 326898 507770 327134
rect 508006 326898 538490 327134
rect 538726 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 31610 295174
rect 31846 294938 62330 295174
rect 62566 294938 93050 295174
rect 93286 294938 123770 295174
rect 124006 294938 154490 295174
rect 154726 294938 185210 295174
rect 185446 294938 215930 295174
rect 216166 294938 246650 295174
rect 246886 294938 277370 295174
rect 277606 294938 308090 295174
rect 308326 294938 338810 295174
rect 339046 294938 369530 295174
rect 369766 294938 400250 295174
rect 400486 294938 430970 295174
rect 431206 294938 461690 295174
rect 461926 294938 492410 295174
rect 492646 294938 523130 295174
rect 523366 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 31610 294854
rect 31846 294618 62330 294854
rect 62566 294618 93050 294854
rect 93286 294618 123770 294854
rect 124006 294618 154490 294854
rect 154726 294618 185210 294854
rect 185446 294618 215930 294854
rect 216166 294618 246650 294854
rect 246886 294618 277370 294854
rect 277606 294618 308090 294854
rect 308326 294618 338810 294854
rect 339046 294618 369530 294854
rect 369766 294618 400250 294854
rect 400486 294618 430970 294854
rect 431206 294618 461690 294854
rect 461926 294618 492410 294854
rect 492646 294618 523130 294854
rect 523366 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 16250 291454
rect 16486 291218 46970 291454
rect 47206 291218 77690 291454
rect 77926 291218 108410 291454
rect 108646 291218 139130 291454
rect 139366 291218 169850 291454
rect 170086 291218 200570 291454
rect 200806 291218 231290 291454
rect 231526 291218 262010 291454
rect 262246 291218 292730 291454
rect 292966 291218 323450 291454
rect 323686 291218 354170 291454
rect 354406 291218 384890 291454
rect 385126 291218 415610 291454
rect 415846 291218 446330 291454
rect 446566 291218 477050 291454
rect 477286 291218 507770 291454
rect 508006 291218 538490 291454
rect 538726 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 16250 291134
rect 16486 290898 46970 291134
rect 47206 290898 77690 291134
rect 77926 290898 108410 291134
rect 108646 290898 139130 291134
rect 139366 290898 169850 291134
rect 170086 290898 200570 291134
rect 200806 290898 231290 291134
rect 231526 290898 262010 291134
rect 262246 290898 292730 291134
rect 292966 290898 323450 291134
rect 323686 290898 354170 291134
rect 354406 290898 384890 291134
rect 385126 290898 415610 291134
rect 415846 290898 446330 291134
rect 446566 290898 477050 291134
rect 477286 290898 507770 291134
rect 508006 290898 538490 291134
rect 538726 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 31610 259174
rect 31846 258938 62330 259174
rect 62566 258938 93050 259174
rect 93286 258938 123770 259174
rect 124006 258938 154490 259174
rect 154726 258938 185210 259174
rect 185446 258938 215930 259174
rect 216166 258938 246650 259174
rect 246886 258938 277370 259174
rect 277606 258938 308090 259174
rect 308326 258938 338810 259174
rect 339046 258938 369530 259174
rect 369766 258938 400250 259174
rect 400486 258938 430970 259174
rect 431206 258938 461690 259174
rect 461926 258938 492410 259174
rect 492646 258938 523130 259174
rect 523366 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 31610 258854
rect 31846 258618 62330 258854
rect 62566 258618 93050 258854
rect 93286 258618 123770 258854
rect 124006 258618 154490 258854
rect 154726 258618 185210 258854
rect 185446 258618 215930 258854
rect 216166 258618 246650 258854
rect 246886 258618 277370 258854
rect 277606 258618 308090 258854
rect 308326 258618 338810 258854
rect 339046 258618 369530 258854
rect 369766 258618 400250 258854
rect 400486 258618 430970 258854
rect 431206 258618 461690 258854
rect 461926 258618 492410 258854
rect 492646 258618 523130 258854
rect 523366 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 16250 255454
rect 16486 255218 46970 255454
rect 47206 255218 77690 255454
rect 77926 255218 108410 255454
rect 108646 255218 139130 255454
rect 139366 255218 169850 255454
rect 170086 255218 200570 255454
rect 200806 255218 231290 255454
rect 231526 255218 262010 255454
rect 262246 255218 292730 255454
rect 292966 255218 323450 255454
rect 323686 255218 354170 255454
rect 354406 255218 384890 255454
rect 385126 255218 415610 255454
rect 415846 255218 446330 255454
rect 446566 255218 477050 255454
rect 477286 255218 507770 255454
rect 508006 255218 538490 255454
rect 538726 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 16250 255134
rect 16486 254898 46970 255134
rect 47206 254898 77690 255134
rect 77926 254898 108410 255134
rect 108646 254898 139130 255134
rect 139366 254898 169850 255134
rect 170086 254898 200570 255134
rect 200806 254898 231290 255134
rect 231526 254898 262010 255134
rect 262246 254898 292730 255134
rect 292966 254898 323450 255134
rect 323686 254898 354170 255134
rect 354406 254898 384890 255134
rect 385126 254898 415610 255134
rect 415846 254898 446330 255134
rect 446566 254898 477050 255134
rect 477286 254898 507770 255134
rect 508006 254898 538490 255134
rect 538726 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 31610 223174
rect 31846 222938 62330 223174
rect 62566 222938 93050 223174
rect 93286 222938 123770 223174
rect 124006 222938 154490 223174
rect 154726 222938 185210 223174
rect 185446 222938 215930 223174
rect 216166 222938 246650 223174
rect 246886 222938 277370 223174
rect 277606 222938 308090 223174
rect 308326 222938 338810 223174
rect 339046 222938 369530 223174
rect 369766 222938 400250 223174
rect 400486 222938 430970 223174
rect 431206 222938 461690 223174
rect 461926 222938 492410 223174
rect 492646 222938 523130 223174
rect 523366 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 31610 222854
rect 31846 222618 62330 222854
rect 62566 222618 93050 222854
rect 93286 222618 123770 222854
rect 124006 222618 154490 222854
rect 154726 222618 185210 222854
rect 185446 222618 215930 222854
rect 216166 222618 246650 222854
rect 246886 222618 277370 222854
rect 277606 222618 308090 222854
rect 308326 222618 338810 222854
rect 339046 222618 369530 222854
rect 369766 222618 400250 222854
rect 400486 222618 430970 222854
rect 431206 222618 461690 222854
rect 461926 222618 492410 222854
rect 492646 222618 523130 222854
rect 523366 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 16250 219454
rect 16486 219218 46970 219454
rect 47206 219218 77690 219454
rect 77926 219218 108410 219454
rect 108646 219218 139130 219454
rect 139366 219218 169850 219454
rect 170086 219218 200570 219454
rect 200806 219218 231290 219454
rect 231526 219218 262010 219454
rect 262246 219218 292730 219454
rect 292966 219218 323450 219454
rect 323686 219218 354170 219454
rect 354406 219218 384890 219454
rect 385126 219218 415610 219454
rect 415846 219218 446330 219454
rect 446566 219218 477050 219454
rect 477286 219218 507770 219454
rect 508006 219218 538490 219454
rect 538726 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 16250 219134
rect 16486 218898 46970 219134
rect 47206 218898 77690 219134
rect 77926 218898 108410 219134
rect 108646 218898 139130 219134
rect 139366 218898 169850 219134
rect 170086 218898 200570 219134
rect 200806 218898 231290 219134
rect 231526 218898 262010 219134
rect 262246 218898 292730 219134
rect 292966 218898 323450 219134
rect 323686 218898 354170 219134
rect 354406 218898 384890 219134
rect 385126 218898 415610 219134
rect 415846 218898 446330 219134
rect 446566 218898 477050 219134
rect 477286 218898 507770 219134
rect 508006 218898 538490 219134
rect 538726 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 31610 187174
rect 31846 186938 62330 187174
rect 62566 186938 93050 187174
rect 93286 186938 123770 187174
rect 124006 186938 154490 187174
rect 154726 186938 185210 187174
rect 185446 186938 215930 187174
rect 216166 186938 246650 187174
rect 246886 186938 277370 187174
rect 277606 186938 308090 187174
rect 308326 186938 338810 187174
rect 339046 186938 369530 187174
rect 369766 186938 400250 187174
rect 400486 186938 430970 187174
rect 431206 186938 461690 187174
rect 461926 186938 492410 187174
rect 492646 186938 523130 187174
rect 523366 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 31610 186854
rect 31846 186618 62330 186854
rect 62566 186618 93050 186854
rect 93286 186618 123770 186854
rect 124006 186618 154490 186854
rect 154726 186618 185210 186854
rect 185446 186618 215930 186854
rect 216166 186618 246650 186854
rect 246886 186618 277370 186854
rect 277606 186618 308090 186854
rect 308326 186618 338810 186854
rect 339046 186618 369530 186854
rect 369766 186618 400250 186854
rect 400486 186618 430970 186854
rect 431206 186618 461690 186854
rect 461926 186618 492410 186854
rect 492646 186618 523130 186854
rect 523366 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 16250 183454
rect 16486 183218 46970 183454
rect 47206 183218 77690 183454
rect 77926 183218 108410 183454
rect 108646 183218 139130 183454
rect 139366 183218 169850 183454
rect 170086 183218 200570 183454
rect 200806 183218 231290 183454
rect 231526 183218 262010 183454
rect 262246 183218 292730 183454
rect 292966 183218 323450 183454
rect 323686 183218 354170 183454
rect 354406 183218 384890 183454
rect 385126 183218 415610 183454
rect 415846 183218 446330 183454
rect 446566 183218 477050 183454
rect 477286 183218 507770 183454
rect 508006 183218 538490 183454
rect 538726 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 16250 183134
rect 16486 182898 46970 183134
rect 47206 182898 77690 183134
rect 77926 182898 108410 183134
rect 108646 182898 139130 183134
rect 139366 182898 169850 183134
rect 170086 182898 200570 183134
rect 200806 182898 231290 183134
rect 231526 182898 262010 183134
rect 262246 182898 292730 183134
rect 292966 182898 323450 183134
rect 323686 182898 354170 183134
rect 354406 182898 384890 183134
rect 385126 182898 415610 183134
rect 415846 182898 446330 183134
rect 446566 182898 477050 183134
rect 477286 182898 507770 183134
rect 508006 182898 538490 183134
rect 538726 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 31610 151174
rect 31846 150938 62330 151174
rect 62566 150938 93050 151174
rect 93286 150938 123770 151174
rect 124006 150938 154490 151174
rect 154726 150938 185210 151174
rect 185446 150938 215930 151174
rect 216166 150938 246650 151174
rect 246886 150938 277370 151174
rect 277606 150938 308090 151174
rect 308326 150938 338810 151174
rect 339046 150938 369530 151174
rect 369766 150938 400250 151174
rect 400486 150938 430970 151174
rect 431206 150938 461690 151174
rect 461926 150938 492410 151174
rect 492646 150938 523130 151174
rect 523366 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 31610 150854
rect 31846 150618 62330 150854
rect 62566 150618 93050 150854
rect 93286 150618 123770 150854
rect 124006 150618 154490 150854
rect 154726 150618 185210 150854
rect 185446 150618 215930 150854
rect 216166 150618 246650 150854
rect 246886 150618 277370 150854
rect 277606 150618 308090 150854
rect 308326 150618 338810 150854
rect 339046 150618 369530 150854
rect 369766 150618 400250 150854
rect 400486 150618 430970 150854
rect 431206 150618 461690 150854
rect 461926 150618 492410 150854
rect 492646 150618 523130 150854
rect 523366 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 16250 147454
rect 16486 147218 46970 147454
rect 47206 147218 77690 147454
rect 77926 147218 108410 147454
rect 108646 147218 139130 147454
rect 139366 147218 169850 147454
rect 170086 147218 200570 147454
rect 200806 147218 231290 147454
rect 231526 147218 262010 147454
rect 262246 147218 292730 147454
rect 292966 147218 323450 147454
rect 323686 147218 354170 147454
rect 354406 147218 384890 147454
rect 385126 147218 415610 147454
rect 415846 147218 446330 147454
rect 446566 147218 477050 147454
rect 477286 147218 507770 147454
rect 508006 147218 538490 147454
rect 538726 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 16250 147134
rect 16486 146898 46970 147134
rect 47206 146898 77690 147134
rect 77926 146898 108410 147134
rect 108646 146898 139130 147134
rect 139366 146898 169850 147134
rect 170086 146898 200570 147134
rect 200806 146898 231290 147134
rect 231526 146898 262010 147134
rect 262246 146898 292730 147134
rect 292966 146898 323450 147134
rect 323686 146898 354170 147134
rect 354406 146898 384890 147134
rect 385126 146898 415610 147134
rect 415846 146898 446330 147134
rect 446566 146898 477050 147134
rect 477286 146898 507770 147134
rect 508006 146898 538490 147134
rect 538726 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 31610 115174
rect 31846 114938 62330 115174
rect 62566 114938 93050 115174
rect 93286 114938 123770 115174
rect 124006 114938 154490 115174
rect 154726 114938 185210 115174
rect 185446 114938 215930 115174
rect 216166 114938 246650 115174
rect 246886 114938 277370 115174
rect 277606 114938 308090 115174
rect 308326 114938 338810 115174
rect 339046 114938 369530 115174
rect 369766 114938 400250 115174
rect 400486 114938 430970 115174
rect 431206 114938 461690 115174
rect 461926 114938 492410 115174
rect 492646 114938 523130 115174
rect 523366 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 31610 114854
rect 31846 114618 62330 114854
rect 62566 114618 93050 114854
rect 93286 114618 123770 114854
rect 124006 114618 154490 114854
rect 154726 114618 185210 114854
rect 185446 114618 215930 114854
rect 216166 114618 246650 114854
rect 246886 114618 277370 114854
rect 277606 114618 308090 114854
rect 308326 114618 338810 114854
rect 339046 114618 369530 114854
rect 369766 114618 400250 114854
rect 400486 114618 430970 114854
rect 431206 114618 461690 114854
rect 461926 114618 492410 114854
rect 492646 114618 523130 114854
rect 523366 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 16250 111454
rect 16486 111218 46970 111454
rect 47206 111218 77690 111454
rect 77926 111218 108410 111454
rect 108646 111218 139130 111454
rect 139366 111218 169850 111454
rect 170086 111218 200570 111454
rect 200806 111218 231290 111454
rect 231526 111218 262010 111454
rect 262246 111218 292730 111454
rect 292966 111218 323450 111454
rect 323686 111218 354170 111454
rect 354406 111218 384890 111454
rect 385126 111218 415610 111454
rect 415846 111218 446330 111454
rect 446566 111218 477050 111454
rect 477286 111218 507770 111454
rect 508006 111218 538490 111454
rect 538726 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 16250 111134
rect 16486 110898 46970 111134
rect 47206 110898 77690 111134
rect 77926 110898 108410 111134
rect 108646 110898 139130 111134
rect 139366 110898 169850 111134
rect 170086 110898 200570 111134
rect 200806 110898 231290 111134
rect 231526 110898 262010 111134
rect 262246 110898 292730 111134
rect 292966 110898 323450 111134
rect 323686 110898 354170 111134
rect 354406 110898 384890 111134
rect 385126 110898 415610 111134
rect 415846 110898 446330 111134
rect 446566 110898 477050 111134
rect 477286 110898 507770 111134
rect 508006 110898 538490 111134
rect 538726 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 31610 79174
rect 31846 78938 62330 79174
rect 62566 78938 93050 79174
rect 93286 78938 123770 79174
rect 124006 78938 154490 79174
rect 154726 78938 185210 79174
rect 185446 78938 215930 79174
rect 216166 78938 246650 79174
rect 246886 78938 277370 79174
rect 277606 78938 308090 79174
rect 308326 78938 338810 79174
rect 339046 78938 369530 79174
rect 369766 78938 400250 79174
rect 400486 78938 430970 79174
rect 431206 78938 461690 79174
rect 461926 78938 492410 79174
rect 492646 78938 523130 79174
rect 523366 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 31610 78854
rect 31846 78618 62330 78854
rect 62566 78618 93050 78854
rect 93286 78618 123770 78854
rect 124006 78618 154490 78854
rect 154726 78618 185210 78854
rect 185446 78618 215930 78854
rect 216166 78618 246650 78854
rect 246886 78618 277370 78854
rect 277606 78618 308090 78854
rect 308326 78618 338810 78854
rect 339046 78618 369530 78854
rect 369766 78618 400250 78854
rect 400486 78618 430970 78854
rect 431206 78618 461690 78854
rect 461926 78618 492410 78854
rect 492646 78618 523130 78854
rect 523366 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 16250 75454
rect 16486 75218 46970 75454
rect 47206 75218 77690 75454
rect 77926 75218 108410 75454
rect 108646 75218 139130 75454
rect 139366 75218 169850 75454
rect 170086 75218 200570 75454
rect 200806 75218 231290 75454
rect 231526 75218 262010 75454
rect 262246 75218 292730 75454
rect 292966 75218 323450 75454
rect 323686 75218 354170 75454
rect 354406 75218 384890 75454
rect 385126 75218 415610 75454
rect 415846 75218 446330 75454
rect 446566 75218 477050 75454
rect 477286 75218 507770 75454
rect 508006 75218 538490 75454
rect 538726 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 16250 75134
rect 16486 74898 46970 75134
rect 47206 74898 77690 75134
rect 77926 74898 108410 75134
rect 108646 74898 139130 75134
rect 139366 74898 169850 75134
rect 170086 74898 200570 75134
rect 200806 74898 231290 75134
rect 231526 74898 262010 75134
rect 262246 74898 292730 75134
rect 292966 74898 323450 75134
rect 323686 74898 354170 75134
rect 354406 74898 384890 75134
rect 385126 74898 415610 75134
rect 415846 74898 446330 75134
rect 446566 74898 477050 75134
rect 477286 74898 507770 75134
rect 508006 74898 538490 75134
rect 538726 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 31610 43174
rect 31846 42938 62330 43174
rect 62566 42938 93050 43174
rect 93286 42938 123770 43174
rect 124006 42938 154490 43174
rect 154726 42938 185210 43174
rect 185446 42938 215930 43174
rect 216166 42938 246650 43174
rect 246886 42938 277370 43174
rect 277606 42938 308090 43174
rect 308326 42938 338810 43174
rect 339046 42938 369530 43174
rect 369766 42938 400250 43174
rect 400486 42938 430970 43174
rect 431206 42938 461690 43174
rect 461926 42938 492410 43174
rect 492646 42938 523130 43174
rect 523366 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 31610 42854
rect 31846 42618 62330 42854
rect 62566 42618 93050 42854
rect 93286 42618 123770 42854
rect 124006 42618 154490 42854
rect 154726 42618 185210 42854
rect 185446 42618 215930 42854
rect 216166 42618 246650 42854
rect 246886 42618 277370 42854
rect 277606 42618 308090 42854
rect 308326 42618 338810 42854
rect 339046 42618 369530 42854
rect 369766 42618 400250 42854
rect 400486 42618 430970 42854
rect 431206 42618 461690 42854
rect 461926 42618 492410 42854
rect 492646 42618 523130 42854
rect 523366 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 16250 39454
rect 16486 39218 46970 39454
rect 47206 39218 77690 39454
rect 77926 39218 108410 39454
rect 108646 39218 139130 39454
rect 139366 39218 169850 39454
rect 170086 39218 200570 39454
rect 200806 39218 231290 39454
rect 231526 39218 262010 39454
rect 262246 39218 292730 39454
rect 292966 39218 323450 39454
rect 323686 39218 354170 39454
rect 354406 39218 384890 39454
rect 385126 39218 415610 39454
rect 415846 39218 446330 39454
rect 446566 39218 477050 39454
rect 477286 39218 507770 39454
rect 508006 39218 538490 39454
rect 538726 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 16250 39134
rect 16486 38898 46970 39134
rect 47206 38898 77690 39134
rect 77926 38898 108410 39134
rect 108646 38898 139130 39134
rect 139366 38898 169850 39134
rect 170086 38898 200570 39134
rect 200806 38898 231290 39134
rect 231526 38898 262010 39134
rect 262246 38898 292730 39134
rect 292966 38898 323450 39134
rect 323686 38898 354170 39134
rect 354406 38898 384890 39134
rect 385126 38898 415610 39134
rect 415846 38898 446330 39134
rect 446566 38898 477050 39134
rect 477286 38898 507770 39134
rect 508006 38898 538490 39134
rect 538726 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use rift2Wrap  i_Rift2Wrap
timestamp 0
transform 1 0 12000 0 1 12000
box 0 0 541520 651526
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 660161 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 660161 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 660161 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 660161 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 660161 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 660161 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 660161 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 660161 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 660161 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 660161 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 660161 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 660161 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 660161 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 660161 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 13103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 660161 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 660161 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 660161 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 660161 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 660161 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 660161 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 660161 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 660161 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 660161 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 660161 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 12068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 663100 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 660161 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 660161 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 12068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 663100 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 660161 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 13103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 660161 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 660161 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 660161 53294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 660161 89294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 660161 125294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 660161 161294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 660161 197294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 660161 233294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 660161 269294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 660161 305294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 660161 341294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 660161 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 660161 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 660161 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 660161 485294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 660161 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 660161 24734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 660161 60734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 660161 96734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 660161 132734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 660161 168734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 660161 204734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 660161 240734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 660161 276734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 660161 312734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 660161 348734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 660161 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 660161 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 660161 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 663100 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 660161 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 660161 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 660161 57014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 663100 93014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 660161 129014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 660161 165014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 663100 201014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 660161 237014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 660161 273014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 663100 309014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 660161 345014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 660161 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 660161 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 660161 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 660161 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 660161 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 660161 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 660161 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 660161 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 660161 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 660161 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 660161 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 660161 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 660161 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 660161 316454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 660161 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 660161 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 660161 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 660161 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 660161 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 660161 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 660161 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 12068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 663100 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 660161 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 660161 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 12068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 663100 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 660161 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 660161 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 660161 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 660161 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 660161 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 660161 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 660161 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 660161 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 660161 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 13103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 660161 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 660161 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 660161 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 660161 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 660161 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 660161 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 660161 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 660161 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 660161 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 660161 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 660161 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 660161 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 660161 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 660161 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 660161 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 660161 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 660161 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 538608 651336 538608 651336 0 vccd1
rlabel metal5 291962 694616 291962 694616 0 vccd2
rlabel metal5 291962 666056 291962 666056 0 vdda1
rlabel metal5 291962 673496 291962 673496 0 vdda2
rlabel metal5 291962 669776 291962 669776 0 vssa1
rlabel metal5 291962 677216 291962 677216 0 vssa2
rlabel via4 523248 655056 523248 655056 0 vssd1
rlabel via4 553424 662496 553424 662496 0 vssd2
rlabel metal2 580198 284869 580198 284869 0 analog_io[0]
rlabel metal2 425148 663476 425148 663476 0 analog_io[10]
rlabel metal2 365026 663476 365026 663476 0 analog_io[11]
rlabel metal2 305134 663476 305134 663476 0 analog_io[12]
rlabel metal2 251482 701940 251482 701940 0 analog_io[13]
rlabel metal2 185456 663476 185456 663476 0 analog_io[14]
rlabel metal2 121486 674155 121486 674155 0 analog_io[15]
rlabel metal2 56626 674461 56626 674461 0 analog_io[16]
rlabel metal3 1878 697340 1878 697340 0 analog_io[17]
rlabel metal3 1878 645116 1878 645116 0 analog_io[18]
rlabel metal3 1878 593028 1878 593028 0 analog_io[19]
rlabel metal2 580198 338351 580198 338351 0 analog_io[1]
rlabel metal3 1924 540804 1924 540804 0 analog_io[20]
rlabel metal3 1924 488716 1924 488716 0 analog_io[21]
rlabel metal3 1878 436628 1878 436628 0 analog_io[22]
rlabel metal3 1878 384404 1878 384404 0 analog_io[23]
rlabel metal3 1878 332316 1878 332316 0 analog_io[24]
rlabel metal3 1924 280092 1924 280092 0 analog_io[25]
rlabel metal3 2200 228004 2200 228004 0 analog_io[26]
rlabel metal3 1832 175916 1832 175916 0 analog_io[27]
rlabel metal3 1878 123692 1878 123692 0 analog_io[28]
rlabel metal2 580198 391153 580198 391153 0 analog_io[2]
rlabel metal2 580198 444601 580198 444601 0 analog_io[3]
rlabel metal2 580198 497403 580198 497403 0 analog_io[4]
rlabel metal2 580198 550885 580198 550885 0 analog_io[5]
rlabel metal2 580198 603653 580198 603653 0 analog_io[6]
rlabel metal3 581908 657356 581908 657356 0 analog_io[7]
rlabel metal2 545162 663476 545162 663476 0 analog_io[8]
rlabel metal2 484994 663476 484994 663476 0 analog_io[9]
rlabel metal2 580198 6715 580198 6715 0 io_in[0]
rlabel metal2 580198 457453 580198 457453 0 io_in[10]
rlabel metal2 580198 510969 580198 510969 0 io_in[11]
rlabel metal2 579830 563703 579830 563703 0 io_in[12]
rlabel metal2 580198 617185 580198 617185 0 io_in[13]
rlabel via2 580198 670701 580198 670701 0 io_in[14]
rlabel metal2 559682 701974 559682 701974 0 io_in[15]
rlabel metal2 469998 663476 469998 663476 0 io_in[16]
rlabel metal2 410060 663476 410060 663476 0 io_in[17]
rlabel metal2 350030 663476 350030 663476 0 io_in[18]
rlabel metal2 290046 663476 290046 663476 0 io_in[19]
rlabel metal2 580198 46597 580198 46597 0 io_in[1]
rlabel metal2 230062 663476 230062 663476 0 io_in[20]
rlabel metal2 170078 663476 170078 663476 0 io_in[21]
rlabel metal2 110140 663476 110140 663476 0 io_in[22]
rlabel metal2 40204 703596 40204 703596 0 io_in[23]
rlabel metal3 1924 684284 1924 684284 0 io_in[24]
rlabel metal3 1924 632060 1924 632060 0 io_in[25]
rlabel metal3 1924 579972 1924 579972 0 io_in[26]
rlabel metal3 1970 527884 1970 527884 0 io_in[27]
rlabel metal3 1970 475660 1970 475660 0 io_in[28]
rlabel metal3 1924 423572 1924 423572 0 io_in[29]
rlabel metal2 580198 86547 580198 86547 0 io_in[2]
rlabel metal3 1878 371348 1878 371348 0 io_in[30]
rlabel metal3 1878 319260 1878 319260 0 io_in[31]
rlabel metal3 1694 267172 1694 267172 0 io_in[32]
rlabel metal3 1740 214948 1740 214948 0 io_in[33]
rlabel metal3 1878 162860 1878 162860 0 io_in[34]
rlabel metal3 1878 110636 1878 110636 0 io_in[35]
rlabel metal3 1878 71604 1878 71604 0 io_in[36]
rlabel metal3 1878 32436 1878 32436 0 io_in[37]
rlabel metal2 580198 126463 580198 126463 0 io_in[3]
rlabel metal2 580198 166073 580198 166073 0 io_in[4]
rlabel via2 580198 205683 580198 205683 0 io_in[5]
rlabel metal2 579830 244919 579830 244919 0 io_in[6]
rlabel metal2 580198 298435 580198 298435 0 io_in[7]
rlabel via2 580198 351917 580198 351917 0 io_in[8]
rlabel metal2 580198 404651 580198 404651 0 io_in[9]
rlabel via2 580198 33099 580198 33099 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal2 580198 537319 580198 537319 0 io_oeb[11]
rlabel metal2 579830 590835 579830 590835 0 io_oeb[12]
rlabel metal2 580198 643569 580198 643569 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal2 499990 663476 499990 663476 0 io_oeb[15]
rlabel metal2 462346 701940 462346 701940 0 io_oeb[16]
rlabel metal2 380022 663476 380022 663476 0 io_oeb[17]
rlabel metal2 332534 701940 332534 701940 0 io_oeb[18]
rlabel metal2 260054 663476 260054 663476 0 io_oeb[19]
rlabel metal2 580198 73049 580198 73049 0 io_oeb[1]
rlabel metal2 200452 663476 200452 663476 0 io_oeb[20]
rlabel metal2 140132 663476 140132 663476 0 io_oeb[21]
rlabel metal2 80194 663476 80194 663476 0 io_oeb[22]
rlabel metal2 20164 663476 20164 663476 0 io_oeb[23]
rlabel metal3 2016 658172 2016 658172 0 io_oeb[24]
rlabel metal3 2016 606084 2016 606084 0 io_oeb[25]
rlabel metal3 1878 553860 1878 553860 0 io_oeb[26]
rlabel metal3 2016 501772 2016 501772 0 io_oeb[27]
rlabel metal3 1924 449548 1924 449548 0 io_oeb[28]
rlabel metal3 1924 397460 1924 397460 0 io_oeb[29]
rlabel metal2 579830 112965 579830 112965 0 io_oeb[2]
rlabel metal3 1878 345372 1878 345372 0 io_oeb[30]
rlabel metal3 1648 293148 1648 293148 0 io_oeb[31]
rlabel metal3 2016 241060 2016 241060 0 io_oeb[32]
rlabel metal3 1878 188836 1878 188836 0 io_oeb[33]
rlabel metal3 1786 136748 1786 136748 0 io_oeb[34]
rlabel metal3 2200 84660 2200 84660 0 io_oeb[35]
rlabel metal3 1556 45492 1556 45492 0 io_oeb[36]
rlabel metal3 1740 6460 1740 6460 0 io_oeb[37]
rlabel metal2 579554 152949 579554 152949 0 io_oeb[3]
rlabel metal2 580198 192185 580198 192185 0 io_oeb[4]
rlabel metal2 580198 232101 580198 232101 0 io_oeb[5]
rlabel metal2 579830 272051 579830 272051 0 io_oeb[6]
rlabel metal2 580198 324785 580198 324785 0 io_oeb[7]
rlabel metal2 580198 378301 580198 378301 0 io_oeb[8]
rlabel metal2 580198 431103 580198 431103 0 io_oeb[9]
rlabel metal2 580014 20213 580014 20213 0 io_out[0]
rlabel metal2 580014 471019 580014 471019 0 io_out[10]
rlabel via2 580198 524467 580198 524467 0 io_out[11]
rlabel metal2 580198 577269 580198 577269 0 io_out[12]
rlabel metal2 580014 630751 580014 630751 0 io_out[13]
rlabel metal2 580198 683519 580198 683519 0 io_out[14]
rlabel metal2 543490 702008 543490 702008 0 io_out[15]
rlabel metal2 455002 663476 455002 663476 0 io_out[16]
rlabel metal2 395018 663476 395018 663476 0 io_out[17]
rlabel metal2 335034 663476 335034 663476 0 io_out[18]
rlabel metal2 275050 663476 275050 663476 0 io_out[19]
rlabel metal2 580198 60163 580198 60163 0 io_out[1]
rlabel metal2 215066 663476 215066 663476 0 io_out[20]
rlabel metal2 155082 663476 155082 663476 0 io_out[21]
rlabel metal2 95282 663476 95282 663476 0 io_out[22]
rlabel metal2 23828 703596 23828 703596 0 io_out[23]
rlabel metal3 1970 671228 1970 671228 0 io_out[24]
rlabel metal3 1970 619140 1970 619140 0 io_out[25]
rlabel metal3 1970 566916 1970 566916 0 io_out[26]
rlabel metal3 1878 514828 1878 514828 0 io_out[27]
rlabel metal3 1878 462604 1878 462604 0 io_out[28]
rlabel metal3 1878 410516 1878 410516 0 io_out[29]
rlabel metal2 580198 100079 580198 100079 0 io_out[2]
rlabel metal3 1648 358428 1648 358428 0 io_out[30]
rlabel metal3 1556 306204 1556 306204 0 io_out[31]
rlabel metal3 1878 254116 1878 254116 0 io_out[32]
rlabel metal3 1878 201892 1878 201892 0 io_out[33]
rlabel metal3 1878 149804 1878 149804 0 io_out[34]
rlabel metal3 2200 97580 2200 97580 0 io_out[35]
rlabel metal3 1740 58548 1740 58548 0 io_out[36]
rlabel metal3 1924 19380 1924 19380 0 io_out[37]
rlabel via2 580198 139349 580198 139349 0 io_out[3]
rlabel metal2 580198 178925 580198 178925 0 io_out[4]
rlabel metal2 580198 218535 580198 218535 0 io_out[5]
rlabel metal2 580198 258485 580198 258485 0 io_out[6]
rlabel metal2 580198 311967 580198 311967 0 io_out[7]
rlabel metal2 580198 364735 580198 364735 0 io_out[8]
rlabel metal2 580198 418217 580198 418217 0 io_out[9]
rlabel metal1 136436 9282 136436 9282 0 la_data_in[0]
rlabel metal2 480562 2642 480562 2642 0 la_data_in[100]
rlabel metal2 484058 3390 484058 3390 0 la_data_in[101]
rlabel metal2 450570 9945 450570 9945 0 la_data_in[102]
rlabel metal2 491142 3356 491142 3356 0 la_data_in[103]
rlabel metal2 456642 9877 456642 9877 0 la_data_in[104]
rlabel metal2 498226 3526 498226 3526 0 la_data_in[105]
rlabel metal1 466486 8228 466486 8228 0 la_data_in[106]
rlabel metal2 505402 3390 505402 3390 0 la_data_in[107]
rlabel metal2 508898 3288 508898 3288 0 la_data_in[108]
rlabel metal2 471822 9843 471822 9843 0 la_data_in[109]
rlabel metal2 161322 2098 161322 2098 0 la_data_in[10]
rlabel metal2 474674 10625 474674 10625 0 la_data_in[110]
rlabel metal2 519570 3492 519570 3492 0 la_data_in[111]
rlabel metal2 523066 2812 523066 2812 0 la_data_in[112]
rlabel metal2 483966 10047 483966 10047 0 la_data_in[113]
rlabel metal2 486236 12036 486236 12036 0 la_data_in[114]
rlabel metal2 488658 6051 488658 6051 0 la_data_in[115]
rlabel metal2 537234 2744 537234 2744 0 la_data_in[116]
rlabel metal2 540822 3458 540822 3458 0 la_data_in[117]
rlabel metal2 544410 4138 544410 4138 0 la_data_in[118]
rlabel metal2 501462 12036 501462 12036 0 la_data_in[119]
rlabel metal1 172592 9486 172592 9486 0 la_data_in[11]
rlabel metal2 505034 9877 505034 9877 0 la_data_in[120]
rlabel metal2 507955 11764 507955 11764 0 la_data_in[121]
rlabel metal2 558578 4104 558578 4104 0 la_data_in[122]
rlabel metal2 562074 2642 562074 2642 0 la_data_in[123]
rlabel metal2 565662 3288 565662 3288 0 la_data_in[124]
rlabel metal2 520214 10761 520214 10761 0 la_data_in[125]
rlabel metal2 523066 9809 523066 9809 0 la_data_in[126]
rlabel metal2 526102 10489 526102 10489 0 la_data_in[127]
rlabel metal2 176640 8364 176640 8364 0 la_data_in[12]
rlabel metal2 171994 1656 171994 1656 0 la_data_in[13]
rlabel metal2 175490 1758 175490 1758 0 la_data_in[14]
rlabel metal2 179078 2132 179078 2132 0 la_data_in[15]
rlabel metal2 182574 1826 182574 1826 0 la_data_in[16]
rlabel metal2 192020 12036 192020 12036 0 la_data_in[17]
rlabel metal2 194918 12036 194918 12036 0 la_data_in[18]
rlabel metal2 193246 1792 193246 1792 0 la_data_in[19]
rlabel metal2 136574 6290 136574 6290 0 la_data_in[1]
rlabel metal2 196834 2064 196834 2064 0 la_data_in[20]
rlabel metal2 200330 1928 200330 1928 0 la_data_in[21]
rlabel metal2 203918 1792 203918 1792 0 la_data_in[22]
rlabel metal2 210082 10251 210082 10251 0 la_data_in[23]
rlabel metal1 212060 9486 212060 9486 0 la_data_in[24]
rlabel metal1 215326 8874 215326 8874 0 la_data_in[25]
rlabel metal2 218086 4342 218086 4342 0 la_data_in[26]
rlabel metal1 221904 9418 221904 9418 0 la_data_in[27]
rlabel metal2 225370 12036 225370 12036 0 la_data_in[28]
rlabel metal2 228521 340 228521 340 0 la_data_in[29]
rlabel metal2 132986 2098 132986 2098 0 la_data_in[2]
rlabel metal1 232024 9486 232024 9486 0 la_data_in[30]
rlabel metal2 235842 1962 235842 1962 0 la_data_in[31]
rlabel metal2 238050 10183 238050 10183 0 la_data_in[32]
rlabel metal2 242926 1911 242926 1911 0 la_data_in[33]
rlabel metal2 246422 1928 246422 1928 0 la_data_in[34]
rlabel metal2 250010 2234 250010 2234 0 la_data_in[35]
rlabel metal2 253506 1928 253506 1928 0 la_data_in[36]
rlabel metal2 257094 1758 257094 1758 0 la_data_in[37]
rlabel metal1 257094 9486 257094 9486 0 la_data_in[38]
rlabel metal2 264178 1996 264178 1996 0 la_data_in[39]
rlabel metal2 136482 2200 136482 2200 0 la_data_in[3]
rlabel metal2 267766 1860 267766 1860 0 la_data_in[40]
rlabel metal2 271262 2064 271262 2064 0 la_data_in[41]
rlabel metal2 274850 1928 274850 1928 0 la_data_in[42]
rlabel metal1 272320 9350 272320 9350 0 la_data_in[43]
rlabel metal1 275172 9418 275172 9418 0 la_data_in[44]
rlabel metal2 277334 10557 277334 10557 0 la_data_in[45]
rlabel metal2 289018 2200 289018 2200 0 la_data_in[46]
rlabel metal2 292606 1962 292606 1962 0 la_data_in[47]
rlabel metal2 296102 1690 296102 1690 0 la_data_in[48]
rlabel metal1 290260 9146 290260 9146 0 la_data_in[49]
rlabel metal2 140070 2030 140070 2030 0 la_data_in[4]
rlabel metal1 293204 9486 293204 9486 0 la_data_in[50]
rlabel metal2 306774 2200 306774 2200 0 la_data_in[51]
rlabel metal2 310270 2234 310270 2234 0 la_data_in[52]
rlabel metal2 313858 1996 313858 1996 0 la_data_in[53]
rlabel metal2 317354 2030 317354 2030 0 la_data_in[54]
rlabel metal1 309810 9520 309810 9520 0 la_data_in[55]
rlabel metal2 310914 10421 310914 10421 0 la_data_in[56]
rlabel metal2 313950 10387 313950 10387 0 la_data_in[57]
rlabel metal2 331423 340 331423 340 0 la_data_in[58]
rlabel metal2 335110 1894 335110 1894 0 la_data_in[59]
rlabel metal2 155434 10693 155434 10693 0 la_data_in[5]
rlabel metal2 338698 1928 338698 1928 0 la_data_in[60]
rlabel metal2 326094 10795 326094 10795 0 la_data_in[61]
rlabel metal2 345782 2098 345782 2098 0 la_data_in[62]
rlabel metal2 349278 1860 349278 1860 0 la_data_in[63]
rlabel metal2 352866 1690 352866 1690 0 la_data_in[64]
rlabel metal2 353418 6018 353418 6018 0 la_data_in[65]
rlabel metal2 341274 10795 341274 10795 0 la_data_in[66]
rlabel metal2 363538 1928 363538 1928 0 la_data_in[67]
rlabel metal2 347346 10659 347346 10659 0 la_data_in[68]
rlabel metal2 370622 1894 370622 1894 0 la_data_in[69]
rlabel metal1 155986 9418 155986 9418 0 la_data_in[6]
rlabel metal2 352038 6527 352038 6527 0 la_data_in[70]
rlabel metal2 356086 10591 356086 10591 0 la_data_in[71]
rlabel metal2 364366 6664 364366 6664 0 la_data_in[72]
rlabel metal2 384790 3288 384790 3288 0 la_data_in[73]
rlabel metal2 370162 8398 370162 8398 0 la_data_in[74]
rlabel metal2 391874 2608 391874 2608 0 la_data_in[75]
rlabel metal2 371450 10625 371450 10625 0 la_data_in[76]
rlabel metal2 398958 3390 398958 3390 0 la_data_in[77]
rlabel metal2 377614 9911 377614 9911 0 la_data_in[78]
rlabel metal2 406042 2574 406042 2574 0 la_data_in[79]
rlabel metal2 157734 6528 157734 6528 0 la_data_in[7]
rlabel metal2 409630 3424 409630 3424 0 la_data_in[80]
rlabel metal2 386446 9843 386446 9843 0 la_data_in[81]
rlabel metal2 389850 10659 389850 10659 0 la_data_in[82]
rlabel metal2 392304 12036 392304 12036 0 la_data_in[83]
rlabel metal2 423798 2608 423798 2608 0 la_data_in[84]
rlabel metal2 427294 4138 427294 4138 0 la_data_in[85]
rlabel metal2 430882 3424 430882 3424 0 la_data_in[86]
rlabel metal1 405720 9486 405720 9486 0 la_data_in[87]
rlabel metal2 407484 12036 407484 12036 0 la_data_in[88]
rlabel metal2 411102 9945 411102 9945 0 la_data_in[89]
rlabel metal2 154238 1996 154238 1996 0 la_data_in[8]
rlabel metal2 445050 2744 445050 2744 0 la_data_in[90]
rlabel metal2 448638 4070 448638 4070 0 la_data_in[91]
rlabel metal2 452134 3322 452134 3322 0 la_data_in[92]
rlabel metal2 422618 12036 422618 12036 0 la_data_in[93]
rlabel metal2 426282 9843 426282 9843 0 la_data_in[94]
rlabel metal2 462806 3254 462806 3254 0 la_data_in[95]
rlabel metal2 466302 2710 466302 2710 0 la_data_in[96]
rlabel metal2 469890 3968 469890 3968 0 la_data_in[97]
rlabel metal2 473478 2676 473478 2676 0 la_data_in[98]
rlabel metal2 476974 3424 476974 3424 0 la_data_in[99]
rlabel metal2 157826 2030 157826 2030 0 la_data_in[9]
rlabel metal1 137632 9486 137632 9486 0 la_data_out[0]
rlabel metal2 481758 2778 481758 2778 0 la_data_out[100]
rlabel metal2 485254 2608 485254 2608 0 la_data_out[101]
rlabel metal2 488842 2676 488842 2676 0 la_data_out[102]
rlabel metal2 467222 7310 467222 7310 0 la_data_out[103]
rlabel metal2 457654 9911 457654 9911 0 la_data_out[104]
rlabel metal2 499422 3322 499422 3322 0 la_data_out[105]
rlabel metal2 503010 2880 503010 2880 0 la_data_out[106]
rlabel metal2 466394 10557 466394 10557 0 la_data_out[107]
rlabel metal2 469430 10285 469430 10285 0 la_data_out[108]
rlabel metal2 513590 3254 513590 3254 0 la_data_out[109]
rlabel metal2 171626 10217 171626 10217 0 la_data_out[10]
rlabel metal2 505034 6153 505034 6153 0 la_data_out[110]
rlabel metal2 520766 3968 520766 3968 0 la_data_out[111]
rlabel metal2 524262 3526 524262 3526 0 la_data_out[112]
rlabel metal2 527850 2846 527850 2846 0 la_data_out[113]
rlabel metal2 488014 10727 488014 10727 0 la_data_out[114]
rlabel metal2 491050 10013 491050 10013 0 la_data_out[115]
rlabel metal2 538430 3424 538430 3424 0 la_data_out[116]
rlabel metal2 542018 2812 542018 2812 0 la_data_out[117]
rlabel metal2 545514 2676 545514 2676 0 la_data_out[118]
rlabel metal2 503194 10625 503194 10625 0 la_data_out[119]
rlabel metal1 173604 8738 173604 8738 0 la_data_out[11]
rlabel metal2 506230 9911 506230 9911 0 la_data_out[120]
rlabel metal2 508500 12036 508500 12036 0 la_data_out[121]
rlabel metal2 559774 2608 559774 2608 0 la_data_out[122]
rlabel metal2 563270 4682 563270 4682 0 la_data_out[123]
rlabel metal2 566858 4002 566858 4002 0 la_data_out[124]
rlabel metal2 520736 12036 520736 12036 0 la_data_out[125]
rlabel metal2 523158 5847 523158 5847 0 la_data_out[126]
rlabel metal2 577438 1928 577438 1928 0 la_data_out[127]
rlabel metal1 176502 9486 176502 9486 0 la_data_out[12]
rlabel metal2 173190 1928 173190 1928 0 la_data_out[13]
rlabel metal2 176686 2098 176686 2098 0 la_data_out[14]
rlabel metal2 180274 1962 180274 1962 0 la_data_out[15]
rlabel metal2 183770 1758 183770 1758 0 la_data_out[16]
rlabel metal2 191958 4963 191958 4963 0 la_data_out[17]
rlabel metal2 190854 1894 190854 1894 0 la_data_out[18]
rlabel metal2 194442 1928 194442 1928 0 la_data_out[19]
rlabel metal2 137126 6018 137126 6018 0 la_data_out[1]
rlabel metal2 197938 2234 197938 2234 0 la_data_out[20]
rlabel metal1 203274 9486 203274 9486 0 la_data_out[21]
rlabel metal1 206586 8738 206586 8738 0 la_data_out[22]
rlabel metal2 211186 10217 211186 10217 0 la_data_out[23]
rlabel metal1 213164 8534 213164 8534 0 la_data_out[24]
rlabel metal1 216430 9486 216430 9486 0 la_data_out[25]
rlabel metal2 219282 5007 219282 5007 0 la_data_out[26]
rlabel metal2 223162 12036 223162 12036 0 la_data_out[27]
rlabel metal2 226474 12036 226474 12036 0 la_data_out[28]
rlabel metal2 229625 340 229625 340 0 la_data_out[29]
rlabel metal2 134182 1656 134182 1656 0 la_data_out[2]
rlabel metal1 233220 9486 233220 9486 0 la_data_out[30]
rlabel metal1 236486 9486 236486 9486 0 la_data_out[31]
rlabel metal2 238694 10251 238694 10251 0 la_data_out[32]
rlabel metal1 243110 8602 243110 8602 0 la_data_out[33]
rlabel metal2 247618 1690 247618 1690 0 la_data_out[34]
rlabel metal2 251206 1826 251206 1826 0 la_data_out[35]
rlabel metal2 254702 1690 254702 1690 0 la_data_out[36]
rlabel metal1 254564 9486 254564 9486 0 la_data_out[37]
rlabel metal2 257278 10285 257278 10285 0 la_data_out[38]
rlabel metal2 265374 1792 265374 1792 0 la_data_out[39]
rlabel metal2 137678 2166 137678 2166 0 la_data_out[3]
rlabel metal2 268870 2098 268870 2098 0 la_data_out[40]
rlabel metal2 272458 1962 272458 1962 0 la_data_out[41]
rlabel metal2 276046 1656 276046 1656 0 la_data_out[42]
rlabel metal1 273470 9282 273470 9282 0 la_data_out[43]
rlabel metal1 276138 9486 276138 9486 0 la_data_out[44]
rlabel metal2 286626 1996 286626 1996 0 la_data_out[45]
rlabel metal2 290214 1928 290214 1928 0 la_data_out[46]
rlabel metal2 293710 2132 293710 2132 0 la_data_out[47]
rlabel metal1 288098 9486 288098 9486 0 la_data_out[48]
rlabel metal1 291594 9350 291594 9350 0 la_data_out[49]
rlabel metal2 141266 2098 141266 2098 0 la_data_out[4]
rlabel metal1 294400 8602 294400 8602 0 la_data_out[50]
rlabel metal2 307970 1894 307970 1894 0 la_data_out[51]
rlabel metal2 311466 2132 311466 2132 0 la_data_out[52]
rlabel metal2 315054 1962 315054 1962 0 la_data_out[53]
rlabel metal2 306406 5950 306406 5950 0 la_data_out[54]
rlabel metal2 308890 10659 308890 10659 0 la_data_out[55]
rlabel metal2 311834 10625 311834 10625 0 la_data_out[56]
rlabel metal2 329222 1724 329222 1724 0 la_data_out[57]
rlabel metal2 332718 1843 332718 1843 0 la_data_out[58]
rlabel metal2 325910 8976 325910 8976 0 la_data_out[59]
rlabel metal2 156446 10591 156446 10591 0 la_data_out[5]
rlabel metal2 330326 5984 330326 5984 0 la_data_out[60]
rlabel metal2 327014 10353 327014 10353 0 la_data_out[61]
rlabel metal2 346978 1996 346978 1996 0 la_data_out[62]
rlabel metal2 350474 1826 350474 1826 0 la_data_out[63]
rlabel metal2 354062 4716 354062 4716 0 la_data_out[64]
rlabel metal2 357558 1928 357558 1928 0 la_data_out[65]
rlabel metal2 361146 1724 361146 1724 0 la_data_out[66]
rlabel metal2 364642 1894 364642 1894 0 la_data_out[67]
rlabel metal2 348358 10693 348358 10693 0 la_data_out[68]
rlabel metal2 371489 340 371489 340 0 la_data_out[69]
rlabel metal1 157412 9078 157412 9078 0 la_data_out[6]
rlabel metal2 354430 10557 354430 10557 0 la_data_out[70]
rlabel metal2 378902 2132 378902 2132 0 la_data_out[71]
rlabel metal2 382398 2030 382398 2030 0 la_data_out[72]
rlabel metal2 385986 2234 385986 2234 0 la_data_out[73]
rlabel metal2 389482 3322 389482 3322 0 la_data_out[74]
rlabel metal2 393070 2948 393070 2948 0 la_data_out[75]
rlabel metal2 371266 5949 371266 5949 0 la_data_out[76]
rlabel metal2 375222 9877 375222 9877 0 la_data_out[77]
rlabel metal2 403650 3356 403650 3356 0 la_data_out[78]
rlabel metal2 407238 1911 407238 1911 0 la_data_out[79]
rlabel metal2 151846 1894 151846 1894 0 la_data_out[7]
rlabel metal2 410826 2642 410826 2642 0 la_data_out[80]
rlabel metal2 386446 6527 386446 6527 0 la_data_out[81]
rlabel metal2 390494 10489 390494 10489 0 la_data_out[82]
rlabel metal2 393714 9809 393714 9809 0 la_data_out[83]
rlabel metal2 424994 3254 424994 3254 0 la_data_out[84]
rlabel metal2 428490 1962 428490 1962 0 la_data_out[85]
rlabel metal2 432078 1707 432078 1707 0 la_data_out[86]
rlabel metal2 405674 10557 405674 10557 0 la_data_out[87]
rlabel metal1 409952 9486 409952 9486 0 la_data_out[88]
rlabel metal2 442658 3356 442658 3356 0 la_data_out[89]
rlabel metal2 155434 1826 155434 1826 0 la_data_out[8]
rlabel metal2 446246 3458 446246 3458 0 la_data_out[90]
rlabel metal2 449834 4036 449834 4036 0 la_data_out[91]
rlabel metal2 420854 10523 420854 10523 0 la_data_out[92]
rlabel metal2 424258 10659 424258 10659 0 la_data_out[93]
rlabel metal2 426758 12036 426758 12036 0 la_data_out[94]
rlabel metal2 464002 1826 464002 1826 0 la_data_out[95]
rlabel metal2 467498 1758 467498 1758 0 la_data_out[96]
rlabel metal2 471086 1996 471086 1996 0 la_data_out[97]
rlabel metal2 474582 1792 474582 1792 0 la_data_out[98]
rlabel metal2 441892 12036 441892 12036 0 la_data_out[99]
rlabel metal2 158930 2064 158930 2064 0 la_data_out[9]
rlabel metal2 133906 6494 133906 6494 0 la_oenb[0]
rlabel metal2 482862 2200 482862 2200 0 la_oenb[100]
rlabel metal2 486450 2166 486450 2166 0 la_oenb[101]
rlabel metal2 489946 2098 489946 2098 0 la_oenb[102]
rlabel metal2 493534 2064 493534 2064 0 la_oenb[103]
rlabel metal2 497122 1843 497122 1843 0 la_oenb[104]
rlabel metal2 500618 2132 500618 2132 0 la_oenb[105]
rlabel metal2 504206 2030 504206 2030 0 la_oenb[106]
rlabel metal2 467774 10523 467774 10523 0 la_oenb[107]
rlabel metal2 469246 5235 469246 5235 0 la_oenb[108]
rlabel metal2 473846 10489 473846 10489 0 la_oenb[109]
rlabel metal2 172638 10659 172638 10659 0 la_oenb[10]
rlabel metal2 518374 1996 518374 1996 0 la_oenb[110]
rlabel metal2 521870 1894 521870 1894 0 la_oenb[111]
rlabel metal2 525458 1928 525458 1928 0 la_oenb[112]
rlabel metal2 485622 10659 485622 10659 0 la_oenb[113]
rlabel metal2 488628 12036 488628 12036 0 la_oenb[114]
rlabel metal2 498226 9486 498226 9486 0 la_oenb[115]
rlabel metal2 539626 1792 539626 1792 0 la_oenb[116]
rlabel metal2 543214 4716 543214 4716 0 la_oenb[117]
rlabel metal2 546710 2234 546710 2234 0 la_oenb[118]
rlabel metal2 504206 10591 504206 10591 0 la_oenb[119]
rlabel metal1 175444 9418 175444 9418 0 la_oenb[11]
rlabel metal2 506752 12036 506752 12036 0 la_oenb[120]
rlabel metal2 557382 1860 557382 1860 0 la_oenb[121]
rlabel metal2 560878 2166 560878 2166 0 la_oenb[122]
rlabel metal2 564466 2132 564466 2132 0 la_oenb[123]
rlabel metal2 518988 12036 518988 12036 0 la_oenb[124]
rlabel metal2 521886 12036 521886 12036 0 la_oenb[125]
rlabel metal2 524784 12036 524784 12036 0 la_oenb[126]
rlabel metal2 578634 1996 578634 1996 0 la_oenb[127]
rlabel metal1 178342 9010 178342 9010 0 la_oenb[12]
rlabel metal2 174294 1826 174294 1826 0 la_oenb[13]
rlabel metal2 177882 1894 177882 1894 0 la_oenb[14]
rlabel metal2 181470 1928 181470 1928 0 la_oenb[15]
rlabel metal2 190824 12036 190824 12036 0 la_oenb[16]
rlabel metal2 193246 5201 193246 5201 0 la_oenb[17]
rlabel metal2 192050 1826 192050 1826 0 la_oenb[18]
rlabel metal2 195638 2166 195638 2166 0 la_oenb[19]
rlabel metal2 138230 6528 138230 6528 0 la_oenb[1]
rlabel metal2 199134 2030 199134 2030 0 la_oenb[20]
rlabel metal2 202722 1826 202722 1826 0 la_oenb[21]
rlabel metal1 207644 9486 207644 9486 0 la_oenb[22]
rlabel metal1 210956 9010 210956 9010 0 la_oenb[23]
rlabel metal1 214360 9486 214360 9486 0 la_oenb[24]
rlabel metal1 217534 9282 217534 9282 0 la_oenb[25]
rlabel metal1 220846 8738 220846 8738 0 la_oenb[26]
rlabel metal2 223783 340 223783 340 0 la_oenb[27]
rlabel metal2 227578 12036 227578 12036 0 la_oenb[28]
rlabel metal2 230858 12036 230858 12036 0 la_oenb[29]
rlabel metal2 135286 2132 135286 2132 0 la_oenb[2]
rlabel metal2 234646 1911 234646 1911 0 la_oenb[30]
rlabel metal1 237544 9418 237544 9418 0 la_oenb[31]
rlabel metal2 241730 1928 241730 1928 0 la_oenb[32]
rlabel metal2 245226 1690 245226 1690 0 la_oenb[33]
rlabel metal2 248623 340 248623 340 0 la_oenb[34]
rlabel metal2 252402 1928 252402 1928 0 la_oenb[35]
rlabel metal2 255898 1996 255898 1996 0 la_oenb[36]
rlabel metal1 255898 8874 255898 8874 0 la_oenb[37]
rlabel metal2 258014 10489 258014 10489 0 la_oenb[38]
rlabel metal2 266570 1928 266570 1928 0 la_oenb[39]
rlabel metal2 138874 2064 138874 2064 0 la_oenb[3]
rlabel metal2 270066 1826 270066 1826 0 la_oenb[40]
rlabel metal2 273654 1996 273654 1996 0 la_oenb[41]
rlabel metal2 277150 1826 277150 1826 0 la_oenb[42]
rlabel metal1 273838 9486 273838 9486 0 la_oenb[43]
rlabel metal2 276506 10285 276506 10285 0 la_oenb[44]
rlabel metal2 287822 2234 287822 2234 0 la_oenb[45]
rlabel metal2 291410 2098 291410 2098 0 la_oenb[46]
rlabel metal2 294906 2030 294906 2030 0 la_oenb[47]
rlabel metal2 288420 9452 288420 9452 0 la_oenb[48]
rlabel metal1 292744 9010 292744 9010 0 la_oenb[49]
rlabel metal2 154606 10489 154606 10489 0 la_oenb[4]
rlabel metal1 295320 9418 295320 9418 0 la_oenb[50]
rlabel metal2 309074 2098 309074 2098 0 la_oenb[51]
rlabel metal2 312662 2064 312662 2064 0 la_oenb[52]
rlabel metal2 303462 10489 303462 10489 0 la_oenb[53]
rlabel metal1 307464 9486 307464 9486 0 la_oenb[54]
rlabel metal2 309902 10795 309902 10795 0 la_oenb[55]
rlabel metal2 312938 10455 312938 10455 0 la_oenb[56]
rlabel metal2 330418 1928 330418 1928 0 la_oenb[57]
rlabel metal2 333914 1962 333914 1962 0 la_oenb[58]
rlabel metal2 337502 1724 337502 1724 0 la_oenb[59]
rlabel metal1 154698 9554 154698 9554 0 la_oenb[5]
rlabel metal2 333270 6154 333270 6154 0 la_oenb[60]
rlabel metal1 331108 9486 331108 9486 0 la_oenb[61]
rlabel metal2 348082 1962 348082 1962 0 la_oenb[62]
rlabel metal2 351670 1962 351670 1962 0 la_oenb[63]
rlabel metal2 353326 6154 353326 6154 0 la_oenb[64]
rlabel metal2 358754 1690 358754 1690 0 la_oenb[65]
rlabel metal2 362342 1962 362342 1962 0 la_oenb[66]
rlabel metal2 346334 10523 346334 10523 0 la_oenb[67]
rlabel metal2 369426 2166 369426 2166 0 la_oenb[68]
rlabel metal2 372922 2098 372922 2098 0 la_oenb[69]
rlabel metal1 158884 9486 158884 9486 0 la_oenb[6]
rlabel metal2 368414 6222 368414 6222 0 la_oenb[70]
rlabel metal2 380006 2064 380006 2064 0 la_oenb[71]
rlabel metal2 361514 10489 361514 10489 0 la_oenb[72]
rlabel metal2 387182 1996 387182 1996 0 la_oenb[73]
rlabel metal2 390678 1962 390678 1962 0 la_oenb[74]
rlabel metal2 370086 12036 370086 12036 0 la_oenb[75]
rlabel metal2 372984 12036 372984 12036 0 la_oenb[76]
rlabel metal1 377200 3978 377200 3978 0 la_oenb[77]
rlabel metal2 404846 1928 404846 1928 0 la_oenb[78]
rlabel metal2 408434 2166 408434 2166 0 la_oenb[79]
rlabel metal2 153042 1928 153042 1928 0 la_oenb[7]
rlabel metal2 411930 2064 411930 2064 0 la_oenb[80]
rlabel metal2 388164 12036 388164 12036 0 la_oenb[81]
rlabel metal2 390586 5507 390586 5507 0 la_oenb[82]
rlabel metal2 422602 1996 422602 1996 0 la_oenb[83]
rlabel metal2 426190 2030 426190 2030 0 la_oenb[84]
rlabel metal2 429686 1894 429686 1894 0 la_oenb[85]
rlabel metal2 403344 12036 403344 12036 0 la_oenb[86]
rlabel metal2 405766 5371 405766 5371 0 la_oenb[87]
rlabel metal2 408526 5201 408526 5201 0 la_oenb[88]
rlabel metal2 443854 2166 443854 2166 0 la_oenb[89]
rlabel metal2 156630 1962 156630 1962 0 la_oenb[8]
rlabel metal2 447442 2064 447442 2064 0 la_oenb[90]
rlabel metal2 450938 4750 450938 4750 0 la_oenb[91]
rlabel metal2 454526 2132 454526 2132 0 la_oenb[92]
rlabel metal2 424902 10557 424902 10557 0 la_oenb[93]
rlabel metal2 461610 2030 461610 2030 0 la_oenb[94]
rlabel metal2 431342 10489 431342 10489 0 la_oenb[95]
rlabel metal2 468694 1962 468694 1962 0 la_oenb[96]
rlabel metal2 472282 1894 472282 1894 0 la_oenb[97]
rlabel metal2 475778 1860 475778 1860 0 la_oenb[98]
rlabel metal2 443088 12036 443088 12036 0 la_oenb[99]
rlabel metal2 160126 1894 160126 1894 0 la_oenb[9]
rlabel metal2 579830 1894 579830 1894 0 user_clock2
rlabel metal2 581026 2030 581026 2030 0 user_irq[0]
rlabel metal2 582222 1843 582222 1843 0 user_irq[1]
rlabel metal2 583418 1962 583418 1962 0 user_irq[2]
rlabel metal2 598 1690 598 1690 0 wb_clk_i
rlabel metal2 1702 2608 1702 2608 0 wb_rst_i
rlabel metal2 2898 1928 2898 1928 0 wbs_ack_o
rlabel metal2 39024 12036 39024 12036 0 wbs_adr_i[0]
rlabel metal2 47886 4070 47886 4070 0 wbs_adr_i[10]
rlabel metal2 76376 12036 76376 12036 0 wbs_adr_i[11]
rlabel metal2 78798 6527 78798 6527 0 wbs_adr_i[12]
rlabel metal2 58466 3968 58466 3968 0 wbs_adr_i[13]
rlabel metal2 62054 2608 62054 2608 0 wbs_adr_i[14]
rlabel metal2 65550 3288 65550 3288 0 wbs_adr_i[15]
rlabel metal2 69138 4002 69138 4002 0 wbs_adr_i[16]
rlabel metal2 94714 10183 94714 10183 0 wbs_adr_i[17]
rlabel metal2 76222 3322 76222 3322 0 wbs_adr_i[18]
rlabel metal2 79718 2574 79718 2574 0 wbs_adr_i[19]
rlabel metal2 43118 12036 43118 12036 0 wbs_adr_i[1]
rlabel metal2 83306 1860 83306 1860 0 wbs_adr_i[20]
rlabel metal2 86894 2166 86894 2166 0 wbs_adr_i[21]
rlabel metal2 90390 2132 90390 2132 0 wbs_adr_i[22]
rlabel metal2 93978 1860 93978 1860 0 wbs_adr_i[23]
rlabel metal2 97474 2064 97474 2064 0 wbs_adr_i[24]
rlabel metal2 119018 12036 119018 12036 0 wbs_adr_i[25]
rlabel metal1 121716 9486 121716 9486 0 wbs_adr_i[26]
rlabel metal2 124338 5439 124338 5439 0 wbs_adr_i[27]
rlabel metal2 111642 1894 111642 1894 0 wbs_adr_i[28]
rlabel metal2 115230 2064 115230 2064 0 wbs_adr_i[29]
rlabel metal2 17066 3968 17066 3968 0 wbs_adr_i[2]
rlabel metal2 118818 1758 118818 1758 0 wbs_adr_i[30]
rlabel metal2 122314 1792 122314 1792 0 wbs_adr_i[31]
rlabel metal2 21850 2642 21850 2642 0 wbs_adr_i[3]
rlabel metal2 55446 12036 55446 12036 0 wbs_adr_i[4]
rlabel metal2 58282 9877 58282 9877 0 wbs_adr_i[5]
rlabel metal2 61196 12036 61196 12036 0 wbs_adr_i[6]
rlabel metal2 37214 3288 37214 3288 0 wbs_adr_i[7]
rlabel metal2 40710 2574 40710 2574 0 wbs_adr_i[8]
rlabel metal2 44298 2064 44298 2064 0 wbs_adr_i[9]
rlabel metal2 4094 1894 4094 1894 0 wbs_cyc_i
rlabel metal2 40312 12036 40312 12036 0 wbs_dat_i[0]
rlabel metal2 74766 12036 74766 12036 0 wbs_dat_i[10]
rlabel metal2 77572 12036 77572 12036 0 wbs_dat_i[11]
rlabel metal2 56074 2200 56074 2200 0 wbs_dat_i[12]
rlabel metal2 59662 1860 59662 1860 0 wbs_dat_i[13]
rlabel metal2 63250 2234 63250 2234 0 wbs_dat_i[14]
rlabel metal2 66746 1894 66746 1894 0 wbs_dat_i[15]
rlabel metal2 70334 1928 70334 1928 0 wbs_dat_i[16]
rlabel metal2 95650 12036 95650 12036 0 wbs_dat_i[17]
rlabel metal2 77418 1826 77418 1826 0 wbs_dat_i[18]
rlabel metal2 80914 1792 80914 1792 0 wbs_dat_i[19]
rlabel metal2 44406 12036 44406 12036 0 wbs_dat_i[1]
rlabel metal2 84502 2030 84502 2030 0 wbs_dat_i[20]
rlabel metal2 87998 2098 87998 2098 0 wbs_dat_i[21]
rlabel metal2 91586 1894 91586 1894 0 wbs_dat_i[22]
rlabel metal2 95174 1758 95174 1758 0 wbs_dat_i[23]
rlabel metal2 98670 1724 98670 1724 0 wbs_dat_i[24]
rlabel metal1 118542 9486 118542 9486 0 wbs_dat_i[25]
rlabel metal2 111918 6154 111918 6154 0 wbs_dat_i[26]
rlabel metal2 109342 2098 109342 2098 0 wbs_dat_i[27]
rlabel metal2 112838 1860 112838 1860 0 wbs_dat_i[28]
rlabel metal2 116426 2234 116426 2234 0 wbs_dat_i[29]
rlabel metal2 18262 2098 18262 2098 0 wbs_dat_i[2]
rlabel metal2 119922 1928 119922 1928 0 wbs_dat_i[30]
rlabel metal2 138230 10625 138230 10625 0 wbs_dat_i[31]
rlabel metal2 23046 4750 23046 4750 0 wbs_dat_i[3]
rlabel metal1 55752 9486 55752 9486 0 wbs_dat_i[4]
rlabel metal2 59386 10693 59386 10693 0 wbs_dat_i[5]
rlabel metal2 62392 12036 62392 12036 0 wbs_dat_i[6]
rlabel metal2 38410 1894 38410 1894 0 wbs_dat_i[7]
rlabel metal2 41906 2132 41906 2132 0 wbs_dat_i[8]
rlabel metal2 45494 1792 45494 1792 0 wbs_dat_i[9]
rlabel metal2 41078 10523 41078 10523 0 wbs_dat_o[0]
rlabel metal2 75486 10489 75486 10489 0 wbs_dat_o[10]
rlabel metal2 78768 12036 78768 12036 0 wbs_dat_o[11]
rlabel metal2 57270 4682 57270 4682 0 wbs_dat_o[12]
rlabel metal2 60858 2166 60858 2166 0 wbs_dat_o[13]
rlabel metal2 64354 4716 64354 4716 0 wbs_dat_o[14]
rlabel metal2 67942 2132 67942 2132 0 wbs_dat_o[15]
rlabel metal2 93994 12036 93994 12036 0 wbs_dat_o[16]
rlabel metal2 75026 2064 75026 2064 0 wbs_dat_o[17]
rlabel metal2 78614 1843 78614 1843 0 wbs_dat_o[18]
rlabel metal2 82110 1758 82110 1758 0 wbs_dat_o[19]
rlabel metal1 44666 9486 44666 9486 0 wbs_dat_o[1]
rlabel metal2 85698 2200 85698 2200 0 wbs_dat_o[20]
rlabel metal2 89194 2234 89194 2234 0 wbs_dat_o[21]
rlabel metal2 92782 4648 92782 4648 0 wbs_dat_o[22]
rlabel metal2 96278 1996 96278 1996 0 wbs_dat_o[23]
rlabel metal2 117990 10523 117990 10523 0 wbs_dat_o[24]
rlabel metal2 121026 10557 121026 10557 0 wbs_dat_o[25]
rlabel metal2 124200 9452 124200 9452 0 wbs_dat_o[26]
rlabel metal2 110538 2132 110538 2132 0 wbs_dat_o[27]
rlabel metal2 114034 2030 114034 2030 0 wbs_dat_o[28]
rlabel metal2 117622 2200 117622 2200 0 wbs_dat_o[29]
rlabel metal2 19458 4784 19458 4784 0 wbs_dat_o[2]
rlabel metal2 121118 1826 121118 1826 0 wbs_dat_o[30]
rlabel metal2 139426 10557 139426 10557 0 wbs_dat_o[31]
rlabel metal2 24242 2200 24242 2200 0 wbs_dat_o[3]
rlabel metal2 57148 12036 57148 12036 0 wbs_dat_o[4]
rlabel metal2 59570 4997 59570 4997 0 wbs_dat_o[5]
rlabel metal2 36018 1928 36018 1928 0 wbs_dat_o[6]
rlabel metal2 39606 1843 39606 1843 0 wbs_dat_o[7]
rlabel metal2 43102 1996 43102 1996 0 wbs_dat_o[8]
rlabel metal2 46690 1962 46690 1962 0 wbs_dat_o[9]
rlabel metal2 41446 5405 41446 5405 0 wbs_sel_i[0]
rlabel metal2 15962 4716 15962 4716 0 wbs_sel_i[1]
rlabel metal2 20654 2030 20654 2030 0 wbs_sel_i[2]
rlabel metal2 25346 4818 25346 4818 0 wbs_sel_i[3]
rlabel metal2 5290 1792 5290 1792 0 wbs_stb_i
rlabel metal2 6486 4648 6486 4648 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
